
`timescale 1ps / 1ps

module jpeg_top_tb;


reg end_of_file_signal;
reg [23:0]data_in;
reg clk;
reg rst;
reg enable;
wire [31:0]JPEG_bitstream;
wire data_ready;
wire [4:0]end_of_file_bitstream_count;
wire eof_data_partial_ready;



// Unit Under Test 
	jpeg_top UUT (
		.end_of_file_signal(end_of_file_signal),
		.data_in(data_in),
		.clk(clk),
		.rst(rst),
		.enable(enable),
		.JPEG_bitstream(JPEG_bitstream),
		.data_ready(data_ready),
		.end_of_file_bitstream_count(end_of_file_bitstream_count),
		.eof_data_partial_ready(eof_data_partial_ready));



initial
begin : STIMUL 
	#0
	rst = 1'b1;
	enable = 1'b0;
	end_of_file_signal = 1'b0;
    #10000; 
	rst = 1'b0;
	enable = 1'b1;
	// data_in holds the red, green, and blue pixel values
	// obtained from the .tif image file

		data_in <= 24'b000100010000010000000110;
#10000;
	data_in <= 24'b000100110000011000001000;
#10000;
	data_in <= 24'b000101100000100100001011;
#10000;
	data_in <= 24'b000101110000101000001100;
#10000;
	data_in <= 24'b000110010000101100001100;
#10000;
	data_in <= 24'b000110000000101000001011;
#10000;
	data_in <= 24'b000110100000101100001001;
#10000;
	data_in <= 24'b000110100000101100001000;
#10000;
	data_in <= 24'b000100100000010100000111;
#10000;
	data_in <= 24'b000100110000011000001000;
#10000;
	data_in <= 24'b000101100000100100001011;
#10000;
	data_in <= 24'b000101110000101000001100;
#10000;
	data_in <= 24'b000110010000101100001100;
#10000;
	data_in <= 24'b000110010000101100001100;
#10000;
	data_in <= 24'b000110110000110000001010;
#10000;
	data_in <= 24'b000110110000110000001001;
#10000;
	data_in <= 24'b000100110000011000001000;
#10000;
	data_in <= 24'b000101000000011100001001;
#10000;
	data_in <= 24'b000101100000100000001001;
#10000;
	data_in <= 24'b000110000000101000001011;
#10000;
	data_in <= 24'b000110000000101000001011;
#10000;
	data_in <= 24'b000110010000101100001100;
#10000;
	data_in <= 24'b000111000000110100001011;
#10000;
	data_in <= 24'b000111010000111000001011;
#10000;
	data_in <= 24'b000100110000011000001000;
#10000;
	data_in <= 24'b000101000000011100001001;
#10000;
	data_in <= 24'b000101100000100000001001;
#10000;
	data_in <= 24'b000101110000100100001010;
#10000;
	data_in <= 24'b000110000000101000001011;
#10000;
	data_in <= 24'b000110010000110000001010;
#10000;
	data_in <= 24'b000111010000111000001011;
#10000;
	data_in <= 24'b000111110001000000001101;
#10000;
	data_in <= 24'b000101010000011100001000;
#10000;
	data_in <= 24'b000101010000011100001000;
#10000;
	data_in <= 24'b000101100000100000001001;
#10000;
	data_in <= 24'b000101110000100100001010;
#10000;
	data_in <= 24'b000110100000101100001001;
#10000;
	data_in <= 24'b000111000000110100001011;
#10000;
	data_in <= 24'b001000000000111100001100;
#10000;
	data_in <= 24'b001000100001000100001110;
#10000;
	data_in <= 24'b000101010000011100001000;
#10000;
	data_in <= 24'b000101100000100000001001;
#10000;
	data_in <= 24'b000101110000100100001010;
#10000;
	data_in <= 24'b000110000000101000001011;
#10000;
	data_in <= 24'b000110110000110000001010;
#10000;
	data_in <= 24'b000111000000110100001011;
#10000;
	data_in <= 24'b001000010001000000001101;
#10000;
	data_in <= 24'b001000100001000100001110;
#10000;
	data_in <= 24'b000101100000100000001001;
#10000;
	data_in <= 24'b000101110000100100001010;
#10000;
	data_in <= 24'b000110100000101100001001;
#10000;
	data_in <= 24'b000110110000110000001010;
#10000;
	data_in <= 24'b000111000000110100001011;
#10000;
	data_in <= 24'b000111010000111000001100;
#10000;
	data_in <= 24'b001000010001000000001101;
#10000;
	data_in <= 24'b001000110001001000001111;
#10000;
	data_in <= 24'b000101110000100100001010;
#10000;
	data_in <= 24'b000110000000101000001011;
#10000;
	data_in <= 24'b000110110000110000001010;
#10000;
	data_in <= 24'b000111000000110100001011;
#10000;
	data_in <= 24'b000111010000111000001100;
#10000;
	data_in <= 24'b000111100000111100001100;
#10000;
	data_in <= 24'b001000100001000100001110;
#10000;
	data_in <= 24'b001000110001001100001101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000111110000111000001011;
#10000;
	data_in <= 24'b000111110000111100001001;
#10000;
	data_in <= 24'b001000110001000100001010;
#10000;
	data_in <= 24'b001001110001010100001110;
#10000;
	data_in <= 24'b001010100001011100001111;
#10000;
	data_in <= 24'b001010110001100000010000;
#10000;
	data_in <= 24'b001011100001100100010001;
#10000;
	data_in <= 24'b001011100001101100010011;
#10000;
	data_in <= 24'b000111100000111000001000;
#10000;
	data_in <= 24'b000111100000111000001000;
#10000;
	data_in <= 24'b001000100001000000001001;
#10000;
	data_in <= 24'b001001110001010100001110;
#10000;
	data_in <= 24'b001010110001100000010000;
#10000;
	data_in <= 24'b001011000001100100010001;
#10000;
	data_in <= 24'b001100000001101100010011;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001000010001000100001011;
#10000;
	data_in <= 24'b001000010001000100001011;
#10000;
	data_in <= 24'b001001000001001000001011;
#10000;
	data_in <= 24'b001001110001010100001110;
#10000;
	data_in <= 24'b001010100001011100001111;
#10000;
	data_in <= 24'b001011000001100100010001;
#10000;
	data_in <= 24'b001011110001101000010010;
#10000;
	data_in <= 24'b001011110001110000010100;
#10000;
	data_in <= 24'b001001000001010000001110;
#10000;
	data_in <= 24'b001000110001001100001101;
#10000;
	data_in <= 24'b001001100001010000001101;
#10000;
	data_in <= 24'b001001110001010100001110;
#10000;
	data_in <= 24'b001010010001011000001110;
#10000;
	data_in <= 24'b001010110001100000010000;
#10000;
	data_in <= 24'b001011100001100100010001;
#10000;
	data_in <= 24'b001011110001101000010010;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001001110001010000001101;
#10000;
	data_in <= 24'b001010000001010100001110;
#10000;
	data_in <= 24'b001010010001011000001110;
#10000;
	data_in <= 24'b001011000001100100010001;
#10000;
	data_in <= 24'b001011110001101100010000;
#10000;
	data_in <= 24'b001100000001110000010001;
#10000;
	data_in <= 24'b001001110001010000001111;
#10000;
	data_in <= 24'b001010000001010100010000;
#10000;
	data_in <= 24'b001010010001011000001111;
#10000;
	data_in <= 24'b001010010001011000001111;
#10000;
	data_in <= 24'b001010100001011100001111;
#10000;
	data_in <= 24'b001011000001100100010001;
#10000;
	data_in <= 24'b001011100001101000001111;
#10000;
	data_in <= 24'b001011100001101000001111;
#10000;
	data_in <= 24'b001010010001011000010001;
#10000;
	data_in <= 24'b001010100001011100010010;
#10000;
	data_in <= 24'b001010110001100000010001;
#10000;
	data_in <= 24'b001010110001100000010001;
#10000;
	data_in <= 24'b001010110001100000010000;
#10000;
	data_in <= 24'b001011000001100100010001;
#10000;
	data_in <= 24'b001011100001101000001111;
#10000;
	data_in <= 24'b001011010001100100001110;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b001010000001011000001111;
#10000;
	data_in <= 24'b001010110001100000010001;
#10000;
	data_in <= 24'b001010110001100000010001;
#10000;
	data_in <= 24'b001011010001101000010010;
#10000;
	data_in <= 24'b001011110001110000010100;
#10000;
	data_in <= 24'b001100010001110100010010;
#10000;
	data_in <= 24'b001100000001110000010001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001100000001110100010101;
#10000;
	data_in <= 24'b001100010010000000010111;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001100100010000000010101;
#10000;
	data_in <= 24'b001100010001111100010100;
#10000;
	data_in <= 24'b001101000010000000010101;
#10000;
	data_in <= 24'b001101010010000100010110;
#10000;
	data_in <= 24'b001100000001110100010101;
#10000;
	data_in <= 24'b001100010010000000010111;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001101000010001000010111;
#10000;
	data_in <= 24'b001100110010000100010110;
#10000;
	data_in <= 24'b001101000010000000010101;
#10000;
	data_in <= 24'b001101000010000000010101;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001100010010000000010111;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001101100010001100011011;
#10000;
	data_in <= 24'b001101110010010100011010;
#10000;
	data_in <= 24'b001101100010010000011001;
#10000;
	data_in <= 24'b001101110010001100011000;
#10000;
	data_in <= 24'b001101100010001000010111;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001100010010000000010111;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001101100010001100011011;
#10000;
	data_in <= 24'b001101110010010100011010;
#10000;
	data_in <= 24'b001110000010011000011011;
#10000;
	data_in <= 24'b001110010010010100011010;
#10000;
	data_in <= 24'b001110010010010100011010;
#10000;
	data_in <= 24'b001100000001111000010011;
#10000;
	data_in <= 24'b001100000001111000010011;
#10000;
	data_in <= 24'b001100010001111100010100;
#10000;
	data_in <= 24'b001100110010000100010110;
#10000;
	data_in <= 24'b001101110010001100011000;
#10000;
	data_in <= 24'b001110010010010100011010;
#10000;
	data_in <= 24'b001111010010011100011100;
#10000;
	data_in <= 24'b001111010010011100011100;
#10000;
	data_in <= 24'b001100000001111000010011;
#10000;
	data_in <= 24'b001100010001111100010100;
#10000;
	data_in <= 24'b001100100010000000010101;
#10000;
	data_in <= 24'b001101000010001000010111;
#10000;
	data_in <= 24'b001110000010010000011001;
#10000;
	data_in <= 24'b001110100010011000011011;
#10000;
	data_in <= 24'b001111100010100000011101;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b001100100001111000010011;
#10000;
	data_in <= 24'b001101000010000000010101;
#10000;
	data_in <= 24'b001101100010001000010111;
#10000;
	data_in <= 24'b001101110010001100011000;
#10000;
	data_in <= 24'b001110000010010000011001;
#10000;
	data_in <= 24'b001110010010010100011010;
#10000;
	data_in <= 24'b001111100010100000011100;
#10000;
	data_in <= 24'b010000000010101000011110;
#10000;
	data_in <= 24'b001100000001110000010001;
#10000;
	data_in <= 24'b001100100001111000010011;
#10000;
	data_in <= 24'b001101010010000100010110;
#10000;
	data_in <= 24'b001101100010001000010111;
#10000;
	data_in <= 24'b001101100010001000010111;
#10000;
	data_in <= 24'b001101100010001000010111;
#10000;
	data_in <= 24'b001110100010010000011000;
#10000;
	data_in <= 24'b001111000010011000011010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001101010001111100010100;
#10000;
	data_in <= 24'b001101010001111100010100;
#10000;
	data_in <= 24'b001101110001111100010011;
#10000;
	data_in <= 24'b001110000010000000010100;
#10000;
	data_in <= 24'b001101110001111100010011;
#10000;
	data_in <= 24'b001101100001111000010010;
#10000;
	data_in <= 24'b001101110001110100010001;
#10000;
	data_in <= 24'b001110000001111000010010;
#10000;
	data_in <= 24'b001101010001111100010100;
#10000;
	data_in <= 24'b001101000001111000010011;
#10000;
	data_in <= 24'b001101110001111100010011;
#10000;
	data_in <= 24'b001110010010000100010101;
#10000;
	data_in <= 24'b001110010010000100010101;
#10000;
	data_in <= 24'b001110000010000000010100;
#10000;
	data_in <= 24'b001110100010000000010100;
#10000;
	data_in <= 24'b001110110010000100010101;
#10000;
	data_in <= 24'b001101100010000000010100;
#10000;
	data_in <= 24'b001101010001111100010011;
#10000;
	data_in <= 24'b001110000010000000010100;
#10000;
	data_in <= 24'b001110100010001000010110;
#10000;
	data_in <= 24'b001110110010001100010111;
#10000;
	data_in <= 24'b001110100010001000010110;
#10000;
	data_in <= 24'b001111000010001000010110;
#10000;
	data_in <= 24'b001111000010001000010110;
#10000;
	data_in <= 24'b001110010010001100010111;
#10000;
	data_in <= 24'b001101110010000100010101;
#10000;
	data_in <= 24'b001110010010000100010101;
#10000;
	data_in <= 24'b001110110010001100010111;
#10000;
	data_in <= 24'b001110110010001100010111;
#10000;
	data_in <= 24'b001110100010001000010110;
#10000;
	data_in <= 24'b001110110010000100010101;
#10000;
	data_in <= 24'b001111000010001000010100;
#10000;
	data_in <= 24'b001110110010010100011001;
#10000;
	data_in <= 24'b001110010010001100010111;
#10000;
	data_in <= 24'b001110100010001000010110;
#10000;
	data_in <= 24'b001110100010001000010110;
#10000;
	data_in <= 24'b001111010010001100010101;
#10000;
	data_in <= 24'b001111000010001000010100;
#10000;
	data_in <= 24'b001111000010001000010100;
#10000;
	data_in <= 24'b001111000010001000010100;
#10000;
	data_in <= 24'b001111010010011100011011;
#10000;
	data_in <= 24'b001110100010010000011000;
#10000;
	data_in <= 24'b001110100010001000010110;
#10000;
	data_in <= 24'b001110110010001100010111;
#10000;
	data_in <= 24'b001111010010001100010101;
#10000;
	data_in <= 24'b001111010010001100010101;
#10000;
	data_in <= 24'b001111100010010000010110;
#10000;
	data_in <= 24'b001111110010010100010111;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010000000010100000011100;
#10000;
	data_in <= 24'b001111010010011000010111;
#10000;
	data_in <= 24'b001111000010010100010110;
#10000;
	data_in <= 24'b001111110010010100010111;
#10000;
	data_in <= 24'b001111110010010100010111;
#10000;
	data_in <= 24'b010000000010011000011000;
#10000;
	data_in <= 24'b010000010010011100011001;
#10000;
	data_in <= 24'b010010010011000100100101;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010000000010100100011010;
#10000;
	data_in <= 24'b001111100010011100011000;
#10000;
	data_in <= 24'b010000000010011000011000;
#10000;
	data_in <= 24'b010000000010011000011000;
#10000;
	data_in <= 24'b010000000010011000011000;
#10000;
	data_in <= 24'b010000010010100000011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001110010001111100010001;
#10000;
	data_in <= 24'b001101010001101100001101;
#10000;
	data_in <= 24'b001110010001111100001111;
#10000;
	data_in <= 24'b001110010001111100001111;
#10000;
	data_in <= 24'b001111000010000000001111;
#10000;
	data_in <= 24'b010000000010010000010011;
#10000;
	data_in <= 24'b001111110010000100001110;
#10000;
	data_in <= 24'b001111000001111000001011;
#10000;
	data_in <= 24'b001111110010010100010111;
#10000;
	data_in <= 24'b001110000001111000010000;
#10000;
	data_in <= 24'b001110010001111100001111;
#10000;
	data_in <= 24'b001101110001110100001101;
#10000;
	data_in <= 24'b001110010001110100001100;
#10000;
	data_in <= 24'b010000000010010000010011;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010001000010011000010011;
#10000;
	data_in <= 24'b001110100010000000010010;
#10000;
	data_in <= 24'b001101110001111000001110;
#10000;
	data_in <= 24'b001111000010001000010010;
#10000;
	data_in <= 24'b001111000010001000010010;
#10000;
	data_in <= 24'b001111100010001000010001;
#10000;
	data_in <= 24'b010000100010011000010101;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b001111010010010000010100;
#10000;
	data_in <= 24'b001101110001111000001110;
#10000;
	data_in <= 24'b001110100010000000010000;
#10000;
	data_in <= 24'b001110010001111100001110;
#10000;
	data_in <= 24'b001110110001111100001110;
#10000;
	data_in <= 24'b010000000010010000010011;
#10000;
	data_in <= 24'b010001000010011000010011;
#10000;
	data_in <= 24'b010001110010100100010110;
#10000;
	data_in <= 24'b001111000010001100010011;
#10000;
	data_in <= 24'b001101100001110100001101;
#10000;
	data_in <= 24'b001110100010000000001111;
#10000;
	data_in <= 24'b001110110010000100010000;
#10000;
	data_in <= 24'b001111000010000000001111;
#10000;
	data_in <= 24'b010000000010010100010001;
#10000;
	data_in <= 24'b010000100010010000010001;
#10000;
	data_in <= 24'b010001010010011100010100;
#10000;
	data_in <= 24'b001110110010001000010010;
#10000;
	data_in <= 24'b001101110001111000001110;
#10000;
	data_in <= 24'b001111100010010000010011;
#10000;
	data_in <= 24'b010000010010011100010110;
#10000;
	data_in <= 24'b010000110010100000010100;
#10000;
	data_in <= 24'b010000110010100000010100;
#10000;
	data_in <= 24'b010000010010001100010000;
#10000;
	data_in <= 24'b010000010010001100010000;
#10000;
	data_in <= 24'b010001000010101100011011;
#10000;
	data_in <= 24'b001111000010010000010010;
#10000;
	data_in <= 24'b001111100010010000010011;
#10000;
	data_in <= 24'b001111100010010000010011;
#10000;
	data_in <= 24'b010000000010010100010001;
#10000;
	data_in <= 24'b010000110010100000010100;
#10000;
	data_in <= 24'b010001000010011000010011;
#10000;
	data_in <= 24'b010001100010100000010101;
#10000;
	data_in <= 24'b010000110010101100011001;
#10000;
	data_in <= 24'b001111000010010000010010;
#10000;
	data_in <= 24'b010000000010011000010101;
#10000;
	data_in <= 24'b010000110010100100011000;
#10000;
	data_in <= 24'b010001010010101000010110;
#10000;
	data_in <= 24'b010001010010101000010110;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010000110010010000001111;
#10000;
	data_in <= 24'b001111110010000000001011;
#10000;
	data_in <= 24'b010001010010011000010001;
#10000;
	data_in <= 24'b010010100010101100010110;
#10000;
	data_in <= 24'b010001100010011100010010;
#10000;
	data_in <= 24'b010010010010101000010101;
#10000;
	data_in <= 24'b010010110010110000010111;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010000110010010000001111;
#10000;
	data_in <= 24'b010000000010000100001100;
#10000;
	data_in <= 24'b010001100010011100010010;
#10000;
	data_in <= 24'b010010010010101000010101;
#10000;
	data_in <= 24'b010001010010011000010001;
#10000;
	data_in <= 24'b010001100010011100010010;
#10000;
	data_in <= 24'b010010010010101000010101;
#10000;
	data_in <= 24'b010000100010010000010001;
#10000;
	data_in <= 24'b010000110010010000001111;
#10000;
	data_in <= 24'b010000010010001000001101;
#10000;
	data_in <= 24'b010001010010011000010001;
#10000;
	data_in <= 24'b010010000010100100010100;
#10000;
	data_in <= 24'b010001000010010100010000;
#10000;
	data_in <= 24'b010001010010011000010001;
#10000;
	data_in <= 24'b010001110010011100010100;
#10000;
	data_in <= 24'b010000100010010000010011;
#10000;
	data_in <= 24'b010000110010010000001111;
#10000;
	data_in <= 24'b010000010010001000001101;
#10000;
	data_in <= 24'b010000110010010000001111;
#10000;
	data_in <= 24'b010001100010011100010010;
#10000;
	data_in <= 24'b010001010010011000010001;
#10000;
	data_in <= 24'b010001100010011100010010;
#10000;
	data_in <= 24'b010010000010100000010101;
#10000;
	data_in <= 24'b010000100010010000010011;
#10000;
	data_in <= 24'b010001100010011000010011;
#10000;
	data_in <= 24'b010000110010001100010000;
#10000;
	data_in <= 24'b010000100010001000001111;
#10000;
	data_in <= 24'b010001000010010000010001;
#10000;
	data_in <= 24'b010001100010011000010011;
#10000;
	data_in <= 24'b010010000010100000010101;
#10000;
	data_in <= 24'b010001110010011100010100;
#10000;
	data_in <= 24'b010000100010010000010011;
#10000;
	data_in <= 24'b010010100010101000010111;
#10000;
	data_in <= 24'b010001110010011100010100;
#10000;
	data_in <= 24'b010001000010010000010001;
#10000;
	data_in <= 24'b010001000010010000010001;
#10000;
	data_in <= 24'b010001100010011000010011;
#10000;
	data_in <= 24'b010001100010011000010011;
#10000;
	data_in <= 24'b010001010010010100010010;
#10000;
	data_in <= 24'b010000010010001100010010;
#10000;
	data_in <= 24'b010010000010101000010111;
#10000;
	data_in <= 24'b010010000010101000010111;
#10000;
	data_in <= 24'b010001110010011100010100;
#10000;
	data_in <= 24'b010001000010010000010001;
#10000;
	data_in <= 24'b010001010010010000010100;
#10000;
	data_in <= 24'b010001000010001100010011;
#10000;
	data_in <= 24'b010000010010001100010010;
#10000;
	data_in <= 24'b010000100010010000010011;
#10000;
	data_in <= 24'b010001100010100000010101;
#10000;
	data_in <= 24'b010010000010101000010111;
#10000;
	data_in <= 24'b010010000010100000010101;
#10000;
	data_in <= 24'b010001010010010100010010;
#10000;
	data_in <= 24'b010001000010001100010011;
#10000;
	data_in <= 24'b010000110010001000010010;
#10000;
	data_in <= 24'b010000010010001100010010;
#10000;
	data_in <= 24'b010000110010011100010110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010001010010011000010111;
#10000;
	data_in <= 24'b010001100010100100011011;
#10000;
	data_in <= 24'b010010010010100000011001;
#10000;
	data_in <= 24'b010010000010011100011000;
#10000;
	data_in <= 24'b010010010010011100010111;
#10000;
	data_in <= 24'b010010010010011100010111;
#10000;
	data_in <= 24'b010001110010011100010100;
#10000;
	data_in <= 24'b010010000010100000010101;
#10000;
	data_in <= 24'b010000110010010000010101;
#10000;
	data_in <= 24'b010001010010100000011010;
#10000;
	data_in <= 24'b010001100010011100011000;
#10000;
	data_in <= 24'b010001110010011000010111;
#10000;
	data_in <= 24'b010010100010100000011000;
#10000;
	data_in <= 24'b010010010010011100010111;
#10000;
	data_in <= 24'b010001010010010100010010;
#10000;
	data_in <= 24'b010001100010011000010011;
#10000;
	data_in <= 24'b010000110010010000010101;
#10000;
	data_in <= 24'b010001010010100000011010;
#10000;
	data_in <= 24'b010010000010100100011010;
#10000;
	data_in <= 24'b010010010010100000011001;
#10000;
	data_in <= 24'b010011000010101000011010;
#10000;
	data_in <= 24'b010010110010100100011001;
#10000;
	data_in <= 24'b010001110010011000010110;
#10000;
	data_in <= 24'b010001100010010100010101;
#10000;
	data_in <= 24'b010000100010010100010110;
#10000;
	data_in <= 24'b010001110010101000011100;
#10000;
	data_in <= 24'b010010010010101000011011;
#10000;
	data_in <= 24'b010010000010100100011010;
#10000;
	data_in <= 24'b010011000010101100011011;
#10000;
	data_in <= 24'b010011100010110000011100;
#10000;
	data_in <= 24'b010010010010100000011000;
#10000;
	data_in <= 24'b010010000010011100010111;
#10000;
	data_in <= 24'b010000110010011000010111;
#10000;
	data_in <= 24'b010001110010101000011100;
#10000;
	data_in <= 24'b010010000010100100011010;
#10000;
	data_in <= 24'b010001100010011100011000;
#10000;
	data_in <= 24'b010010100010100100011010;
#10000;
	data_in <= 24'b010011000010101100011100;
#10000;
	data_in <= 24'b010010110010101000011010;
#10000;
	data_in <= 24'b010010010010100000011000;
#10000;
	data_in <= 24'b010000110010011000010111;
#10000;
	data_in <= 24'b010001100010101100011101;
#10000;
	data_in <= 24'b010010100010101100011100;
#10000;
	data_in <= 24'b010001100010011100011000;
#10000;
	data_in <= 24'b010010100010100100011010;
#10000;
	data_in <= 24'b010011010010110000011101;
#10000;
	data_in <= 24'b010011010010110000011100;
#10000;
	data_in <= 24'b010011000010101100011011;
#10000;
	data_in <= 24'b010000110010011000010111;
#10000;
	data_in <= 24'b010001110010110100011101;
#10000;
	data_in <= 24'b010010110010110000011101;
#10000;
	data_in <= 24'b010001110010100000011001;
#10000;
	data_in <= 24'b010010100010100100011010;
#10000;
	data_in <= 24'b010011100010101100011101;
#10000;
	data_in <= 24'b010011100010110100011110;
#10000;
	data_in <= 24'b010011100010110100011110;
#10000;
	data_in <= 24'b010000000010001100010100;
#10000;
	data_in <= 24'b010001100010110000011100;
#10000;
	data_in <= 24'b010010110010110000011101;
#10000;
	data_in <= 24'b010001100010011100011000;
#10000;
	data_in <= 24'b010010010010011000011000;
#10000;
	data_in <= 24'b010011000010100100011011;
#10000;
	data_in <= 24'b010011000010101100011100;
#10000;
	data_in <= 24'b010011010010110000011101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010001110010100100010110;
#10000;
	data_in <= 24'b010000100010010000010001;
#10000;
	data_in <= 24'b010000100010010000010001;
#10000;
	data_in <= 24'b010001010010011100010100;
#10000;
	data_in <= 24'b010001100010010100010101;
#10000;
	data_in <= 24'b010000110010001000010010;
#10000;
	data_in <= 24'b010010000010001100010101;
#10000;
	data_in <= 24'b010011000010100100011011;
#10000;
	data_in <= 24'b010001010010011100010100;
#10000;
	data_in <= 24'b010000100010010000010001;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010001010010011100010100;
#10000;
	data_in <= 24'b010001100010010100010101;
#10000;
	data_in <= 24'b010000110010001000010010;
#10000;
	data_in <= 24'b010001010010001000010100;
#10000;
	data_in <= 24'b010010000010010100010111;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010000100010011000010101;
#10000;
	data_in <= 24'b010001100010100000010111;
#10000;
	data_in <= 24'b010010000010011100010111;
#10000;
	data_in <= 24'b010001100010010100010101;
#10000;
	data_in <= 24'b010001100010001100010101;
#10000;
	data_in <= 24'b010001100010010100010110;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010001000010011000010011;
#10000;
	data_in <= 24'b010001000010100000010111;
#10000;
	data_in <= 24'b010001010010100100011000;
#10000;
	data_in <= 24'b010001110010100100011000;
#10000;
	data_in <= 24'b010010010010100000011000;
#10000;
	data_in <= 24'b010010100010011100011001;
#10000;
	data_in <= 24'b010010000010011100010111;
#10000;
	data_in <= 24'b010001000010011000010101;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010001000010100000010111;
#10000;
	data_in <= 24'b010000110010011100010110;
#10000;
	data_in <= 24'b010001100010100000010111;
#10000;
	data_in <= 24'b010010010010100000011000;
#10000;
	data_in <= 24'b010010010010011000011000;
#10000;
	data_in <= 24'b010001110010011000010110;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010000110010011100010110;
#10000;
	data_in <= 24'b010000100010011000010101;
#10000;
	data_in <= 24'b010001000010011000010101;
#10000;
	data_in <= 24'b010001000010011000010101;
#10000;
	data_in <= 24'b010001100010010100010110;
#10000;
	data_in <= 24'b010001000010001100010011;
#10000;
	data_in <= 24'b010001100010100000010111;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010000100010011000010101;
#10000;
	data_in <= 24'b010000110010011100010110;
#10000;
	data_in <= 24'b010001100010100000010111;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010001100010010100010101;
#10000;
	data_in <= 24'b010001100010010100010101;
#10000;
	data_in <= 24'b010010000010011100010111;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010001100010101000011001;
#10000;
	data_in <= 24'b010010100010110000011011;
#10000;
	data_in <= 24'b010010010010101100011010;
#10000;
	data_in <= 24'b010010100010100100011001;
#10000;
	data_in <= 24'b010010100010100100011001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001111110010000100010000;
#10000;
	data_in <= 24'b010000000010001100010100;
#10000;
	data_in <= 24'b010000100010001000010111;
#10000;
	data_in <= 24'b001111110001111100011001;
#10000;
	data_in <= 24'b010000010010001100100010;
#10000;
	data_in <= 24'b010000110010101100101101;
#10000;
	data_in <= 24'b001111110010101000101101;
#10000;
	data_in <= 24'b001101010010010000101000;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010001010010100000011001;
#10000;
	data_in <= 24'b010001010010010100011010;
#10000;
	data_in <= 24'b010000000010000000011011;
#10000;
	data_in <= 24'b010000100010010000100011;
#10000;
	data_in <= 24'b010001010010101000101101;
#10000;
	data_in <= 24'b001111110010100100101110;
#10000;
	data_in <= 24'b001101110010001100101000;
#10000;
	data_in <= 24'b010000110010011100010110;
#10000;
	data_in <= 24'b010000010010011100010111;
#10000;
	data_in <= 24'b010000100010010000011001;
#10000;
	data_in <= 24'b001111110010000100011100;
#10000;
	data_in <= 24'b010000110010010000100111;
#10000;
	data_in <= 24'b010001110010101100110001;
#10000;
	data_in <= 24'b010001000010110000110100;
#10000;
	data_in <= 24'b001111110010100000110000;
#10000;
	data_in <= 24'b001111110010001100010010;
#10000;
	data_in <= 24'b001111100010010000010011;
#10000;
	data_in <= 24'b010000000010000100011000;
#10000;
	data_in <= 24'b001111110010000000011101;
#10000;
	data_in <= 24'b010001000010010100101000;
#10000;
	data_in <= 24'b010010100010101100110100;
#10000;
	data_in <= 24'b010010010010111000111000;
#10000;
	data_in <= 24'b010001010010110000110110;
#10000;
	data_in <= 24'b010000110010011100010110;
#10000;
	data_in <= 24'b010000010010011100010110;
#10000;
	data_in <= 24'b010000100010010100011100;
#10000;
	data_in <= 24'b010000110010010000100001;
#10000;
	data_in <= 24'b010001100010011100101010;
#10000;
	data_in <= 24'b010010100010101100110100;
#10000;
	data_in <= 24'b010011000010101100111001;
#10000;
	data_in <= 24'b010010000010110000111001;
#10000;
	data_in <= 24'b010001100010101000011001;
#10000;
	data_in <= 24'b010001010010101100011010;
#10000;
	data_in <= 24'b010001100010101000011111;
#10000;
	data_in <= 24'b010001100010100000100011;
#10000;
	data_in <= 24'b010010000010100100101010;
#10000;
	data_in <= 24'b010011000010101100110010;
#10000;
	data_in <= 24'b010100010010111000111100;
#10000;
	data_in <= 24'b010100000011000101000000;
#10000;
	data_in <= 24'b010010000010101000011001;
#10000;
	data_in <= 24'b010001110010101100011010;
#10000;
	data_in <= 24'b010001100010101100011101;
#10000;
	data_in <= 24'b010001100010100100100000;
#10000;
	data_in <= 24'b010001110010100000100101;
#10000;
	data_in <= 24'b010010110010101100110000;
#10000;
	data_in <= 24'b010100110011000100111100;
#10000;
	data_in <= 24'b010101010011011001000101;
#10000;
	data_in <= 24'b010010110010101000011011;
#10000;
	data_in <= 24'b010010010010101000011011;
#10000;
	data_in <= 24'b010001110010101000011011;
#10000;
	data_in <= 24'b010001000010100100011011;
#10000;
	data_in <= 24'b010000110010011000011111;
#10000;
	data_in <= 24'b010010000010100100101000;
#10000;
	data_in <= 24'b010100010011000000110111;
#10000;
	data_in <= 24'b010101100011011101000110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001110100010010100101000;
#10000;
	data_in <= 24'b001111100010010100101001;
#10000;
	data_in <= 24'b001111000001110100100000;
#10000;
	data_in <= 24'b010000100001111100100011;
#10000;
	data_in <= 24'b010000110010000100100010;
#10000;
	data_in <= 24'b010000000010000100100010;
#10000;
	data_in <= 24'b001100100001101000011010;
#10000;
	data_in <= 24'b001101010010000000011111;
#10000;
	data_in <= 24'b001101010001111100100100;
#10000;
	data_in <= 24'b001110100010001100100111;
#10000;
	data_in <= 24'b010001010010011000101001;
#10000;
	data_in <= 24'b010001100010010100101001;
#10000;
	data_in <= 24'b001110110001101100011100;
#10000;
	data_in <= 24'b010000100010001100100100;
#10000;
	data_in <= 24'b001111010010010100100101;
#10000;
	data_in <= 24'b001101010010000000011111;
#10000;
	data_in <= 24'b001101110010000100100110;
#10000;
	data_in <= 24'b010000010010101000101110;
#10000;
	data_in <= 24'b001111010010001000100101;
#10000;
	data_in <= 24'b001110110001111100011111;
#10000;
	data_in <= 24'b010000000010000100100010;
#10000;
	data_in <= 24'b010001110010101100101011;
#10000;
	data_in <= 24'b010000000010010100101000;
#10000;
	data_in <= 24'b001111110010011100100111;
#10000;
	data_in <= 24'b001111100010011100101111;
#10000;
	data_in <= 24'b010001000010111000110011;
#10000;
	data_in <= 24'b001110000010000100100101;
#10000;
	data_in <= 24'b001110010010001100100101;
#10000;
	data_in <= 24'b010001010010110100101111;
#10000;
	data_in <= 24'b010010100010111100110010;
#10000;
	data_in <= 24'b010000000010010100101001;
#10000;
	data_in <= 24'b010010010010111000110001;
#10000;
	data_in <= 24'b010000100010101000110110;
#10000;
	data_in <= 24'b001111110010101000110011;
#10000;
	data_in <= 24'b010000000010111000110101;
#10000;
	data_in <= 24'b010001110011011000111010;
#10000;
	data_in <= 24'b010000100010111000110011;
#10000;
	data_in <= 24'b010001110011000000110101;
#10000;
	data_in <= 24'b010010100010111000110100;
#10000;
	data_in <= 24'b010010110010110100110010;
#10000;
	data_in <= 24'b010001110010110100111101;
#10000;
	data_in <= 24'b010000100011000000111101;
#10000;
	data_in <= 24'b001111100011001000111110;
#10000;
	data_in <= 24'b010000010011011001000000;
#10000;
	data_in <= 24'b001111110011000100111100;
#10000;
	data_in <= 24'b010010100011011001000010;
#10000;
	data_in <= 24'b010011000011001100111101;
#10000;
	data_in <= 24'b010010110010111100110101;
#10000;
	data_in <= 24'b010010110011001001000110;
#10000;
	data_in <= 24'b010001010011010001001001;
#10000;
	data_in <= 24'b001110110011001001000111;
#10000;
	data_in <= 24'b010000010011101101001110;
#10000;
	data_in <= 24'b010001110011111101010000;
#10000;
	data_in <= 24'b010011100100000101010001;
#10000;
	data_in <= 24'b010011000011010101000100;
#10000;
	data_in <= 24'b010011010011010000111110;
#10000;
	data_in <= 24'b010011000011010001001100;
#10000;
	data_in <= 24'b001110100010101101000111;
#10000;
	data_in <= 24'b010000100011110101011010;
#10000;
	data_in <= 24'b010110000101010001110001;
#10000;
	data_in <= 24'b010011000100100001100001;
#10000;
	data_in <= 24'b010011000100001101011000;
#10000;
	data_in <= 24'b010100000011110101010000;
#10000;
	data_in <= 24'b010011100011011001000010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001110000010000000100000;
#10000;
	data_in <= 24'b001110100010000000100000;
#10000;
	data_in <= 24'b001110100010000000100000;
#10000;
	data_in <= 24'b001110100010000000100000;
#10000;
	data_in <= 24'b001111010010000100100000;
#10000;
	data_in <= 24'b001111010010000100100000;
#10000;
	data_in <= 24'b001111000010000000011111;
#10000;
	data_in <= 24'b001110110001111100011110;
#10000;
	data_in <= 24'b001111000010010000100100;
#10000;
	data_in <= 24'b001111010010010000100010;
#10000;
	data_in <= 24'b001111010010001100100011;
#10000;
	data_in <= 24'b001111010010010000100010;
#10000;
	data_in <= 24'b010000000010010000100011;
#10000;
	data_in <= 24'b010000000010010100100001;
#10000;
	data_in <= 24'b001111110010001100100010;
#10000;
	data_in <= 24'b001111100010001100011111;
#10000;
	data_in <= 24'b010000000010011100100101;
#10000;
	data_in <= 24'b001111110010011000100010;
#10000;
	data_in <= 24'b001111100010010100100011;
#10000;
	data_in <= 24'b001111100010010100100001;
#10000;
	data_in <= 24'b010000010010011000100010;
#10000;
	data_in <= 24'b010000000010011000100000;
#10000;
	data_in <= 24'b001111110010010000100000;
#10000;
	data_in <= 24'b001111110010010100011111;
#10000;
	data_in <= 24'b010000010010100000100110;
#10000;
	data_in <= 24'b010000000010011100100011;
#10000;
	data_in <= 24'b001111110010011000100010;
#10000;
	data_in <= 24'b001111110010011100100001;
#10000;
	data_in <= 24'b010000010010011100100001;
#10000;
	data_in <= 24'b010000000010011000100000;
#10000;
	data_in <= 24'b001111110010010100011111;
#10000;
	data_in <= 24'b001111100010010000011101;
#10000;
	data_in <= 24'b010000110010101000101000;
#10000;
	data_in <= 24'b010000100010101000100100;
#10000;
	data_in <= 24'b010000010010100100100011;
#10000;
	data_in <= 24'b010000010010100100100011;
#10000;
	data_in <= 24'b010000100010100000100010;
#10000;
	data_in <= 24'b010000100010100000100001;
#10000;
	data_in <= 24'b010000000010011000011111;
#10000;
	data_in <= 24'b010000000010011100011101;
#10000;
	data_in <= 24'b010001000010101100101001;
#10000;
	data_in <= 24'b010000110010101100100101;
#10000;
	data_in <= 24'b010000100010101000100100;
#10000;
	data_in <= 24'b010000010010100100100011;
#10000;
	data_in <= 24'b010000110010100100100011;
#10000;
	data_in <= 24'b010000100010100000100001;
#10000;
	data_in <= 24'b010000010010100000011110;
#10000;
	data_in <= 24'b010000000010011100011101;
#10000;
	data_in <= 24'b010001000010100100101100;
#10000;
	data_in <= 24'b010000110010101000100110;
#10000;
	data_in <= 24'b010000010010100000100100;
#10000;
	data_in <= 24'b010000000010100000100010;
#10000;
	data_in <= 24'b010000100010100000100010;
#10000;
	data_in <= 24'b010000010010011100100000;
#10000;
	data_in <= 24'b010000100010011100011101;
#10000;
	data_in <= 24'b010000100010011100011101;
#10000;
	data_in <= 24'b010000110010101000101110;
#10000;
	data_in <= 24'b010000110010101000101000;
#10000;
	data_in <= 24'b010000100010100100100111;
#10000;
	data_in <= 24'b010000010010100000100100;
#10000;
	data_in <= 24'b010000100010011100100011;
#10000;
	data_in <= 24'b010000100010100000100010;
#10000;
	data_in <= 24'b010000110010011100100000;
#10000;
	data_in <= 24'b010000100010011100011101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001110000001110100011001;
#10000;
	data_in <= 24'b001110100001111100011011;
#10000;
	data_in <= 24'b001110010010000000011110;
#10000;
	data_in <= 24'b001101110001111000011100;
#10000;
	data_in <= 24'b001100110001110000011010;
#10000;
	data_in <= 24'b001101000001110100011011;
#10000;
	data_in <= 24'b001101010001111000011100;
#10000;
	data_in <= 24'b001101010001111000011100;
#10000;
	data_in <= 24'b001111000010000100011101;
#10000;
	data_in <= 24'b001111000010000100011101;
#10000;
	data_in <= 24'b001110010010000000011100;
#10000;
	data_in <= 24'b001101100001110100011001;
#10000;
	data_in <= 24'b001100100001101100011001;
#10000;
	data_in <= 24'b001100110001110100011000;
#10000;
	data_in <= 24'b001101000001110100011011;
#10000;
	data_in <= 24'b001101010001111100011010;
#10000;
	data_in <= 24'b001111010010001100011101;
#10000;
	data_in <= 24'b001111000010001000011100;
#10000;
	data_in <= 24'b001110000010000000011010;
#10000;
	data_in <= 24'b001101100001111000011000;
#10000;
	data_in <= 24'b001101100001110100011001;
#10000;
	data_in <= 24'b001101110001111100011001;
#10000;
	data_in <= 24'b001101010001111100011010;
#10000;
	data_in <= 24'b001101000001111000011000;
#10000;
	data_in <= 24'b001110110010000100011011;
#10000;
	data_in <= 24'b001110110010000100011010;
#10000;
	data_in <= 24'b001110000010000000011010;
#10000;
	data_in <= 24'b001110000010000000011010;
#10000;
	data_in <= 24'b001110100010001000011100;
#10000;
	data_in <= 24'b001110100010001000011100;
#10000;
	data_in <= 24'b001110000010000000011010;
#10000;
	data_in <= 24'b001100100001110000010110;
#10000;
	data_in <= 24'b001111000010001000011011;
#10000;
	data_in <= 24'b001110110010001000011000;
#10000;
	data_in <= 24'b001110100010000000011001;
#10000;
	data_in <= 24'b001110110010000100011010;
#10000;
	data_in <= 24'b001111010010001100011100;
#10000;
	data_in <= 24'b001110110010010000011100;
#10000;
	data_in <= 24'b001110000010000100011001;
#10000;
	data_in <= 24'b001101000001110100010101;
#10000;
	data_in <= 24'b001111110010011000011100;
#10000;
	data_in <= 24'b001111010010010000011010;
#10000;
	data_in <= 24'b001110110010001000011000;
#10000;
	data_in <= 24'b001110100010000100010111;
#10000;
	data_in <= 24'b001110110010000100011010;
#10000;
	data_in <= 24'b001111000010001000011011;
#10000;
	data_in <= 24'b001110010001111100011000;
#10000;
	data_in <= 24'b001101000001110100010101;
#10000;
	data_in <= 24'b010000000010010100011011;
#10000;
	data_in <= 24'b001111110010010000011010;
#10000;
	data_in <= 24'b001111010010001000011000;
#10000;
	data_in <= 24'b001111000010000100010111;
#10000;
	data_in <= 24'b001111010010001000011000;
#10000;
	data_in <= 24'b001111000010001100011001;
#10000;
	data_in <= 24'b001110010001111100011000;
#10000;
	data_in <= 24'b001101010001101100010100;
#10000;
	data_in <= 24'b001111010010001000011000;
#10000;
	data_in <= 24'b001111010010001000011000;
#10000;
	data_in <= 24'b001111100010001100011001;
#10000;
	data_in <= 24'b001111100010001100011001;
#10000;
	data_in <= 24'b010000000010010100011011;
#10000;
	data_in <= 24'b001111110010010000011010;
#10000;
	data_in <= 24'b001110110001111100011000;
#10000;
	data_in <= 24'b001101010001101100010100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000110100000101100001001;
#10000;
	data_in <= 24'b000110110000110000001010;
#10000;
	data_in <= 24'b000111000000110100001011;
#10000;
	data_in <= 24'b000111000000110100001011;
#10000;
	data_in <= 24'b000111110000111000001011;
#10000;
	data_in <= 24'b001000000000111100001100;
#10000;
	data_in <= 24'b001001000001000100001110;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b000110110000110000001010;
#10000;
	data_in <= 24'b000111000000110100001011;
#10000;
	data_in <= 24'b000111010000111000001100;
#10000;
	data_in <= 24'b000111010000111000001100;
#10000;
	data_in <= 24'b001000000000111100001100;
#10000;
	data_in <= 24'b001000100001000100001110;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b001001110001010000001111;
#10000;
	data_in <= 24'b000111100000110100001010;
#10000;
	data_in <= 24'b000111100000110100001010;
#10000;
	data_in <= 24'b001000000000111100001100;
#10000;
	data_in <= 24'b001000010001000000001101;
#10000;
	data_in <= 24'b001000100001000100001110;
#10000;
	data_in <= 24'b001001000001001100010000;
#10000;
	data_in <= 24'b001010000001010100010000;
#10000;
	data_in <= 24'b001010100001011100010010;
#10000;
	data_in <= 24'b000111100000110100001010;
#10000;
	data_in <= 24'b000111110000111000001011;
#10000;
	data_in <= 24'b001000000000111100001100;
#10000;
	data_in <= 24'b001000010001000000001101;
#10000;
	data_in <= 24'b001000110001001000001111;
#10000;
	data_in <= 24'b001001010001010100001111;
#10000;
	data_in <= 24'b001010010001011000010001;
#10000;
	data_in <= 24'b001010110001100000010011;
#10000;
	data_in <= 24'b000111010000110000001001;
#10000;
	data_in <= 24'b000111100000110100001010;
#10000;
	data_in <= 24'b001000000000111100001100;
#10000;
	data_in <= 24'b001000010001000000001101;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001001110001010000001111;
#10000;
	data_in <= 24'b001010100001011100010010;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b000111010000110000001001;
#10000;
	data_in <= 24'b000111100000110100001010;
#10000;
	data_in <= 24'b001000000000111100001100;
#10000;
	data_in <= 24'b001000100001000100001110;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b001010000001010100010000;
#10000;
	data_in <= 24'b001010110001100100010010;
#10000;
	data_in <= 24'b001011010001101100010100;
#10000;
	data_in <= 24'b000111100000110100001010;
#10000;
	data_in <= 24'b000111110000111000001011;
#10000;
	data_in <= 24'b001000110001000000001011;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001001110001010000001111;
#10000;
	data_in <= 24'b001010010001011000010001;
#10000;
	data_in <= 24'b001011010001101000010011;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b000111110000111000001011;
#10000;
	data_in <= 24'b001000000000111100001100;
#10000;
	data_in <= 24'b001001000001000100001100;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b001001110001010000001111;
#10000;
	data_in <= 24'b001010100001011100010010;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001001110001010100001110;
#10000;
	data_in <= 24'b001010110001100000010001;
#10000;
	data_in <= 24'b001011010001101000010010;
#10000;
	data_in <= 24'b001100010001110000010100;
#10000;
	data_in <= 24'b001100010001110000010100;
#10000;
	data_in <= 24'b001100000001110000010001;
#10000;
	data_in <= 24'b001011110001101100010000;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b001100000001110100010101;
#10000;
	data_in <= 24'b001100000001110100010101;
#10000;
	data_in <= 24'b001100010001110000010100;
#10000;
	data_in <= 24'b001100010001110000010100;
#10000;
	data_in <= 24'b001100100001111000010011;
#10000;
	data_in <= 24'b001101000010000000010101;
#10000;
	data_in <= 24'b001011000001100100010010;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100100001111100010111;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001100000001110000010001;
#10000;
	data_in <= 24'b001100000001110000010001;
#10000;
	data_in <= 24'b001101000010000000010101;
#10000;
	data_in <= 24'b001110010010010100011010;
#10000;
	data_in <= 24'b001010110001100000010001;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001100000001110100010101;
#10000;
	data_in <= 24'b001100010001110100010010;
#10000;
	data_in <= 24'b001100100001111000010011;
#10000;
	data_in <= 24'b001101100010001000010111;
#10000;
	data_in <= 24'b001110110010011100011100;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100100001111100010111;
#10000;
	data_in <= 24'b001100110010000000011000;
#10000;
	data_in <= 24'b001101010010000100010110;
#10000;
	data_in <= 24'b001101100010001000010111;
#10000;
	data_in <= 24'b001110000010010000011001;
#10000;
	data_in <= 24'b001110100010011000011011;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001100110010000000011000;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001110000010010000011001;
#10000;
	data_in <= 24'b001110010010010100011010;
#10000;
	data_in <= 24'b001110000010010000011001;
#10000;
	data_in <= 24'b001110000010010000011001;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001100100001111100010111;
#10000;
	data_in <= 24'b001101100010000100011001;
#10000;
	data_in <= 24'b001110000010001100011011;
#10000;
	data_in <= 24'b001110010010010100011010;
#10000;
	data_in <= 24'b001110010010010100011010;
#10000;
	data_in <= 24'b001110000010010000011001;
#10000;
	data_in <= 24'b001101110010001100011000;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001100110010000000011000;
#10000;
	data_in <= 24'b001110000010001100011011;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011100011100;
#10000;
	data_in <= 24'b001110110010011100011100;
#10000;
	data_in <= 24'b001110110010011100011100;
#10000;
	data_in <= 24'b001110110010011100011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001100110001111100010100;
#10000;
	data_in <= 24'b001100010001110100010010;
#10000;
	data_in <= 24'b001101000001111000010010;
#10000;
	data_in <= 24'b001101110010000100010101;
#10000;
	data_in <= 24'b001110010010001100010111;
#10000;
	data_in <= 24'b001110000010001000010110;
#10000;
	data_in <= 24'b001110100010010000011000;
#10000;
	data_in <= 24'b001111000010011000011010;
#10000;
	data_in <= 24'b001101000010000000010101;
#10000;
	data_in <= 24'b001100110001111100010100;
#10000;
	data_in <= 24'b001101100010000000010100;
#10000;
	data_in <= 24'b001110000010001000010110;
#10000;
	data_in <= 24'b001110010010001100010111;
#10000;
	data_in <= 24'b001110100010010000011000;
#10000;
	data_in <= 24'b001110110010010100011001;
#10000;
	data_in <= 24'b001111000010011000011010;
#10000;
	data_in <= 24'b001101110010000100010101;
#10000;
	data_in <= 24'b001110000010001000010110;
#10000;
	data_in <= 24'b001110010010001100010111;
#10000;
	data_in <= 24'b001110000010001000010110;
#10000;
	data_in <= 24'b001110010010001100010111;
#10000;
	data_in <= 24'b001110110010010100011001;
#10000;
	data_in <= 24'b001111100010011100011000;
#10000;
	data_in <= 24'b001111100010011100011000;
#10000;
	data_in <= 24'b001110000010001000010110;
#10000;
	data_in <= 24'b001110100010010000011000;
#10000;
	data_in <= 24'b001110110010010100011001;
#10000;
	data_in <= 24'b001110010010001100010111;
#10000;
	data_in <= 24'b001110100010010000011000;
#10000;
	data_in <= 24'b001111000010011000011010;
#10000;
	data_in <= 24'b001111110010100000011001;
#10000;
	data_in <= 24'b001111100010011100011000;
#10000;
	data_in <= 24'b001110010010001100010111;
#10000;
	data_in <= 24'b001110110010010100011001;
#10000;
	data_in <= 24'b001111010010010100011001;
#10000;
	data_in <= 24'b001111000010010000011000;
#10000;
	data_in <= 24'b001111000010010100010110;
#10000;
	data_in <= 24'b001111110010100000011001;
#10000;
	data_in <= 24'b010000000010100100011010;
#10000;
	data_in <= 24'b001111100010011100011000;
#10000;
	data_in <= 24'b001110100010010000011000;
#10000;
	data_in <= 24'b001110110010010100011001;
#10000;
	data_in <= 24'b001111010010010100011001;
#10000;
	data_in <= 24'b001111010010010100011001;
#10000;
	data_in <= 24'b001111100010011100011000;
#10000;
	data_in <= 24'b001111110010100000011001;
#10000;
	data_in <= 24'b010000000010100100011010;
#10000;
	data_in <= 24'b010000000010100100011010;
#10000;
	data_in <= 24'b001110110010010100011001;
#10000;
	data_in <= 24'b001111010010010100011001;
#10000;
	data_in <= 24'b001111010010010100011001;
#10000;
	data_in <= 24'b001111110010011100011011;
#10000;
	data_in <= 24'b001111110010100000011001;
#10000;
	data_in <= 24'b010000000010100100011010;
#10000;
	data_in <= 24'b010000010010101000011011;
#10000;
	data_in <= 24'b010000100010101100011100;
#10000;
	data_in <= 24'b001111000010011000011011;
#10000;
	data_in <= 24'b001111000010010000011000;
#10000;
	data_in <= 24'b001111010010010100011001;
#10000;
	data_in <= 24'b010000000010100000011100;
#10000;
	data_in <= 24'b010000010010100100011101;
#10000;
	data_in <= 24'b010000000010100100011010;
#10000;
	data_in <= 24'b010000010010101000011011;
#10000;
	data_in <= 24'b010001000010110100011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010000110010110000011101;
#10000;
	data_in <= 24'b010001000010110100011110;
#10000;
	data_in <= 24'b010001000010101000011100;
#10000;
	data_in <= 24'b010000100010100000011010;
#10000;
	data_in <= 24'b010001000010101000011100;
#10000;
	data_in <= 24'b010000110010100100011011;
#10000;
	data_in <= 24'b010000110010101000011010;
#10000;
	data_in <= 24'b010001100010110100011101;
#10000;
	data_in <= 24'b001111110010100000011001;
#10000;
	data_in <= 24'b010000110010110000011101;
#10000;
	data_in <= 24'b010010000010111000100000;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010001110010110100011111;
#10000;
	data_in <= 24'b010001010010110000011100;
#10000;
	data_in <= 24'b010001100010110100011101;
#10000;
	data_in <= 24'b001111110010100000011001;
#10000;
	data_in <= 24'b010000110010110000011101;
#10000;
	data_in <= 24'b010001100010110000011110;
#10000;
	data_in <= 24'b010001110010110100011111;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010001110010111000011110;
#10000;
	data_in <= 24'b010001110010111000011110;
#10000;
	data_in <= 24'b010010010011000000100000;
#10000;
	data_in <= 24'b010000010010101000011011;
#10000;
	data_in <= 24'b010000110010110000011101;
#10000;
	data_in <= 24'b010001000010101000011100;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010001110010111000011110;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010000110010100100011011;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010001100010110100011101;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010001100010110000011110;
#10000;
	data_in <= 24'b010001110010110100011111;
#10000;
	data_in <= 24'b010001100010110100011101;
#10000;
	data_in <= 24'b010001110010111000011110;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010010010011000000100000;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010001110010110100011111;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010010011000000100000;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010011100011010100100101;
#10000;
	data_in <= 24'b010001000010101000011100;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010011110011011000100110;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010011010011010000100100;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010011110011011000100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010001010010110100011011;
#10000;
	data_in <= 24'b010001110010111100011101;
#10000;
	data_in <= 24'b010001010010101100011010;
#10000;
	data_in <= 24'b010001010010101100011010;
#10000;
	data_in <= 24'b010011000011000100011101;
#10000;
	data_in <= 24'b010010010010111000011010;
#10000;
	data_in <= 24'b010001010010011100010100;
#10000;
	data_in <= 24'b010010000010101000010111;
#10000;
	data_in <= 24'b010010010011000100011111;
#10000;
	data_in <= 24'b010010010011000100011111;
#10000;
	data_in <= 24'b010001110010110100011100;
#10000;
	data_in <= 24'b010001110010110100011100;
#10000;
	data_in <= 24'b010011000011000100011101;
#10000;
	data_in <= 24'b010010010010111000011010;
#10000;
	data_in <= 24'b010010000010101000010111;
#10000;
	data_in <= 24'b010010110010110100011010;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010010010010111100011110;
#10000;
	data_in <= 24'b010010000010111000011101;
#10000;
	data_in <= 24'b010010110011000000011100;
#10000;
	data_in <= 24'b010010100010111100011011;
#10000;
	data_in <= 24'b010010000010110100011001;
#10000;
	data_in <= 24'b010010110011000000011100;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010100011000000011111;
#10000;
	data_in <= 24'b010010010010111100011110;
#10000;
	data_in <= 24'b010010110010111100011110;
#10000;
	data_in <= 24'b010010100010111100011011;
#10000;
	data_in <= 24'b010010110011000000011100;
#10000;
	data_in <= 24'b010011000011000100011101;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010110011000100100001;
#10000;
	data_in <= 24'b010010110011000100100000;
#10000;
	data_in <= 24'b010011000011000000011111;
#10000;
	data_in <= 24'b010011000011000000011111;
#10000;
	data_in <= 24'b010011010011001000011110;
#10000;
	data_in <= 24'b010011010011001000011110;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011100011001000100001;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010100000011010100100001;
#10000;
	data_in <= 24'b010011010011001000011110;
#10000;
	data_in <= 24'b010011100011010000100110;
#10000;
	data_in <= 24'b010010110011000100100011;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011100011001000100001;
#10000;
	data_in <= 24'b010100000011010000100011;
#10000;
	data_in <= 24'b010100010011011000100010;
#10000;
	data_in <= 24'b010011000011000100011101;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011010011000100100000;
#10000;
	data_in <= 24'b010100000011010000100011;
#10000;
	data_in <= 24'b010100010011011000100010;
#10000;
	data_in <= 24'b010010110011000000011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010001100010100000010101;
#10000;
	data_in <= 24'b010010000010101000010111;
#10000;
	data_in <= 24'b010001110010100100010110;
#10000;
	data_in <= 24'b010001000010011000010011;
#10000;
	data_in <= 24'b010001100010100000010111;
#10000;
	data_in <= 24'b010010010010101100011010;
#10000;
	data_in <= 24'b010001100010100000010111;
#10000;
	data_in <= 24'b001111100010001000010001;
#10000;
	data_in <= 24'b010010110010110100011010;
#10000;
	data_in <= 24'b010011100011000000011101;
#10000;
	data_in <= 24'b010011010010111100011100;
#10000;
	data_in <= 24'b010010000010101000010111;
#10000;
	data_in <= 24'b010001100010100000010111;
#10000;
	data_in <= 24'b010001110010100100011000;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b001111110010001100010010;
#10000;
	data_in <= 24'b010010110010110100011010;
#10000;
	data_in <= 24'b010100000011001000011111;
#10000;
	data_in <= 24'b010100010011001100100000;
#10000;
	data_in <= 24'b010010110010110100011010;
#10000;
	data_in <= 24'b010001110010100100010110;
#10000;
	data_in <= 24'b010001100010100000010101;
#10000;
	data_in <= 24'b010001000010100100010101;
#10000;
	data_in <= 24'b010000110010100000010100;
#10000;
	data_in <= 24'b010010110010110100011010;
#10000;
	data_in <= 24'b010100100011010000100001;
#10000;
	data_in <= 24'b010101010011011100100100;
#10000;
	data_in <= 24'b010100000011001000011111;
#10000;
	data_in <= 24'b010010100010110000011001;
#10000;
	data_in <= 24'b010010000010101000010111;
#10000;
	data_in <= 24'b010001110010110000011000;
#10000;
	data_in <= 24'b010001110010110000011000;
#10000;
	data_in <= 24'b010011100011000100011100;
#10000;
	data_in <= 24'b010101010011100000100011;
#10000;
	data_in <= 24'b010110010011110000100111;
#10000;
	data_in <= 24'b010101010011100000100011;
#10000;
	data_in <= 24'b010011010011001000011101;
#10000;
	data_in <= 24'b010010010010111000011001;
#10000;
	data_in <= 24'b010010000010110100011001;
#10000;
	data_in <= 24'b010010000010110100011001;
#10000;
	data_in <= 24'b010011000010111100011010;
#10000;
	data_in <= 24'b010100010011010000011111;
#10000;
	data_in <= 24'b010101010011100000100011;
#10000;
	data_in <= 24'b010101000011011100100010;
#10000;
	data_in <= 24'b010011100011001100011110;
#10000;
	data_in <= 24'b010011000011000100011100;
#10000;
	data_in <= 24'b010010100010111100011011;
#10000;
	data_in <= 24'b010010010010111000011010;
#10000;
	data_in <= 24'b010010100010110100011000;
#10000;
	data_in <= 24'b010011000010111100011010;
#10000;
	data_in <= 24'b010011000011000100011100;
#10000;
	data_in <= 24'b010011010011001000011101;
#10000;
	data_in <= 24'b010011010011001000011101;
#10000;
	data_in <= 24'b010011010011001000011101;
#10000;
	data_in <= 24'b010010110011000000011011;
#10000;
	data_in <= 24'b010010010010111000011001;
#10000;
	data_in <= 24'b010011100011000000011101;
#10000;
	data_in <= 24'b010011010011000000011011;
#10000;
	data_in <= 24'b010010100010111100011011;
#10000;
	data_in <= 24'b010010100010111100011010;
#10000;
	data_in <= 24'b010011000011000100011101;
#10000;
	data_in <= 24'b010011000011000100011100;
#10000;
	data_in <= 24'b010010010010111000011010;
#10000;
	data_in <= 24'b010010000010101100010110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010010000010101100011100;
#10000;
	data_in <= 24'b010001010010101100011011;
#10000;
	data_in <= 24'b010010110010110000011101;
#10000;
	data_in <= 24'b010010000010100100011010;
#10000;
	data_in <= 24'b010011110010110000011110;
#10000;
	data_in <= 24'b010010100010011100011001;
#10000;
	data_in <= 24'b010011010010101100011011;
#10000;
	data_in <= 24'b010100000010111100011111;
#10000;
	data_in <= 24'b010001100010101000011001;
#10000;
	data_in <= 24'b010001100010100100011010;
#10000;
	data_in <= 24'b010010100010101100011100;
#10000;
	data_in <= 24'b010010010010100000011001;
#10000;
	data_in <= 24'b010100010010111000100000;
#10000;
	data_in <= 24'b010011010010101000011100;
#10000;
	data_in <= 24'b010011010010101100011011;
#10000;
	data_in <= 24'b010011000010101000011010;
#10000;
	data_in <= 24'b010000100010011100010011;
#10000;
	data_in <= 24'b010001010010100100011000;
#10000;
	data_in <= 24'b010010100010110000011011;
#10000;
	data_in <= 24'b010010100010100100011001;
#10000;
	data_in <= 24'b010100110011000100100001;
#10000;
	data_in <= 24'b010100110010111100011111;
#10000;
	data_in <= 24'b010100110010111100011111;
#10000;
	data_in <= 24'b010011110010110100011101;
#10000;
	data_in <= 24'b010000110010100000010100;
#10000;
	data_in <= 24'b010001110010100100010110;
#10000;
	data_in <= 24'b010011100010110100011101;
#10000;
	data_in <= 24'b010011100010110000011100;
#10000;
	data_in <= 24'b010101110011001100100011;
#10000;
	data_in <= 24'b010100100010111000011110;
#10000;
	data_in <= 24'b010101000011000000100000;
#10000;
	data_in <= 24'b010101010011000100100001;
#10000;
	data_in <= 24'b010010000010110100011000;
#10000;
	data_in <= 24'b010010000010101100010110;
#10000;
	data_in <= 24'b010011010010110100011010;
#10000;
	data_in <= 24'b010100010011000000011101;
#10000;
	data_in <= 24'b010110110011011100100101;
#10000;
	data_in <= 24'b010101100011000000011110;
#10000;
	data_in <= 24'b010101000010111000011100;
#10000;
	data_in <= 24'b010100100010111000011100;
#10000;
	data_in <= 24'b010010100010111100011010;
#10000;
	data_in <= 24'b010001100010100100010100;
#10000;
	data_in <= 24'b010010100010101000010111;
#10000;
	data_in <= 24'b010100110010111100011101;
#10000;
	data_in <= 24'b011001000011111000101100;
#10000;
	data_in <= 24'b010111110011100100100111;
#10000;
	data_in <= 24'b010110010011001100100001;
#10000;
	data_in <= 24'b010100110010110100011011;
#10000;
	data_in <= 24'b010010010010110000010111;
#10000;
	data_in <= 24'b010001110010101000010101;
#10000;
	data_in <= 24'b010010010010101000010101;
#10000;
	data_in <= 24'b010011100010101100010111;
#10000;
	data_in <= 24'b011000000011101000101000;
#10000;
	data_in <= 24'b011001000011110000101010;
#10000;
	data_in <= 24'b011000010011100100100111;
#10000;
	data_in <= 24'b010101110011000100011111;
#10000;
	data_in <= 24'b010001110010101000010101;
#10000;
	data_in <= 24'b010011000010110100011000;
#10000;
	data_in <= 24'b010011000010110100011000;
#10000;
	data_in <= 24'b010001100010010100010001;
#10000;
	data_in <= 24'b010101000010111000011100;
#10000;
	data_in <= 24'b010110100011010000100010;
#10000;
	data_in <= 24'b010111010011011100100101;
#10000;
	data_in <= 24'b010101110011000100011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010010010010100000011000;
#10000;
	data_in <= 24'b010001010010011100010110;
#10000;
	data_in <= 24'b010001100010100000010111;
#10000;
	data_in <= 24'b010010000010101000011001;
#10000;
	data_in <= 24'b010010110010101000011010;
#10000;
	data_in <= 24'b010010110010101000011010;
#10000;
	data_in <= 24'b010011000010101000011010;
#10000;
	data_in <= 24'b010011100010101100011101;
#10000;
	data_in <= 24'b010011000010101000011010;
#10000;
	data_in <= 24'b010011000010101100011011;
#10000;
	data_in <= 24'b010010110010101000011010;
#10000;
	data_in <= 24'b010010000010101000011001;
#10000;
	data_in <= 24'b010011000010101100011011;
#10000;
	data_in <= 24'b010011110010111000011110;
#10000;
	data_in <= 24'b010100000010111000011110;
#10000;
	data_in <= 24'b010011010010101100011011;
#10000;
	data_in <= 24'b010011100010110000011100;
#10000;
	data_in <= 24'b010011110010111000011110;
#10000;
	data_in <= 24'b010011100010111000011011;
#10000;
	data_in <= 24'b010010110010101100011000;
#10000;
	data_in <= 24'b010011010010110100011010;
#10000;
	data_in <= 24'b010100010011000100011110;
#10000;
	data_in <= 24'b010100100011000100011110;
#10000;
	data_in <= 24'b010011010010101100011011;
#10000;
	data_in <= 24'b010100010010110100011101;
#10000;
	data_in <= 24'b010100010010111100011111;
#10000;
	data_in <= 24'b010100000010111100011100;
#10000;
	data_in <= 24'b010011000010110000011001;
#10000;
	data_in <= 24'b010011000010110000011001;
#10000;
	data_in <= 24'b010011110011000000011011;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010011010010110000011001;
#10000;
	data_in <= 24'b010100010010110100011011;
#10000;
	data_in <= 24'b010011110010111000011011;
#10000;
	data_in <= 24'b010011110010111000011011;
#10000;
	data_in <= 24'b010011110010111000011011;
#10000;
	data_in <= 24'b010011010010110000011000;
#10000;
	data_in <= 24'b010011000010101100010111;
#10000;
	data_in <= 24'b010100000010110100011001;
#10000;
	data_in <= 24'b010100100010111100011011;
#10000;
	data_in <= 24'b010101010010111100011101;
#10000;
	data_in <= 24'b010100010010110100011011;
#10000;
	data_in <= 24'b010011110010111000011011;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010011110010111000011010;
#10000;
	data_in <= 24'b010011010010110000011000;
#10000;
	data_in <= 24'b010100000010111000010111;
#10000;
	data_in <= 24'b010100110011000000011100;
#10000;
	data_in <= 24'b010101100011000000011110;
#10000;
	data_in <= 24'b010100110010111100011101;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010011110010111000011010;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010100010011000100011010;
#10000;
	data_in <= 24'b010100110011000100011010;
#10000;
	data_in <= 24'b010100010011000100011010;
#10000;
	data_in <= 24'b010101100011000000011110;
#10000;
	data_in <= 24'b010101000011000000011110;
#10000;
	data_in <= 24'b010100100010111100011011;
#10000;
	data_in <= 24'b010011010010110000011000;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010101010011010100011110;
#10000;
	data_in <= 24'b010101100011001100011111;
#10000;
	data_in <= 24'b010011110010111100011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100010010111000100001;
#10000;
	data_in <= 24'b010010010010011100011010;
#10000;
	data_in <= 24'b010001110010100100011000;
#10000;
	data_in <= 24'b010010110010111100011110;
#10000;
	data_in <= 24'b010010110010111000011111;
#10000;
	data_in <= 24'b010001100010100100100010;
#10000;
	data_in <= 24'b010011100010111100110010;
#10000;
	data_in <= 24'b010110010011101001001001;
#10000;
	data_in <= 24'b010100010010111000100001;
#10000;
	data_in <= 24'b010011100010101100011110;
#10000;
	data_in <= 24'b010011000010101100011011;
#10000;
	data_in <= 24'b010011000010111000011011;
#10000;
	data_in <= 24'b010010110010110100011010;
#10000;
	data_in <= 24'b010010000010101100011101;
#10000;
	data_in <= 24'b010010100010110000101011;
#10000;
	data_in <= 24'b010011010011001000111100;
#10000;
	data_in <= 24'b010100000010101000011110;
#10000;
	data_in <= 24'b010011110010110000011111;
#10000;
	data_in <= 24'b010011100010111000011011;
#10000;
	data_in <= 24'b010010100010110100011000;
#10000;
	data_in <= 24'b010010100010110100011000;
#10000;
	data_in <= 24'b010010110010111100011110;
#10000;
	data_in <= 24'b010010110010111000101001;
#10000;
	data_in <= 24'b010001110010110100110011;
#10000;
	data_in <= 24'b010100000010101100011101;
#10000;
	data_in <= 24'b010011110010110000011110;
#10000;
	data_in <= 24'b010011110010111000011011;
#10000;
	data_in <= 24'b010011010010111000010111;
#10000;
	data_in <= 24'b010011000011000000011000;
#10000;
	data_in <= 24'b010011100011001000100001;
#10000;
	data_in <= 24'b010011010011001000101000;
#10000;
	data_in <= 24'b010010000011000000110010;
#10000;
	data_in <= 24'b010100010010111100011111;
#10000;
	data_in <= 24'b010011110010110100011101;
#10000;
	data_in <= 24'b010011110010111000011011;
#10000;
	data_in <= 24'b010011110011000000011011;
#10000;
	data_in <= 24'b010011100011000100011100;
#10000;
	data_in <= 24'b010011010011000100100000;
#10000;
	data_in <= 24'b010010110011001100100111;
#10000;
	data_in <= 24'b010010010011001100101110;
#10000;
	data_in <= 24'b010100000010111100011100;
#10000;
	data_in <= 24'b010011010010110000011001;
#10000;
	data_in <= 24'b010011010010110000011001;
#10000;
	data_in <= 24'b010100010011000000011101;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010011010011000000100001;
#10000;
	data_in <= 24'b010011000011010000101000;
#10000;
	data_in <= 24'b010011110011100000110000;
#10000;
	data_in <= 24'b010011010010111000011001;
#10000;
	data_in <= 24'b010011000010110100011000;
#10000;
	data_in <= 24'b010011100010110100011010;
#10000;
	data_in <= 24'b010100100011000000100000;
#10000;
	data_in <= 24'b010100110011001000100011;
#10000;
	data_in <= 24'b010011110011001000100100;
#10000;
	data_in <= 24'b010011100011011000101010;
#10000;
	data_in <= 24'b010100000011101000101111;
#10000;
	data_in <= 24'b010011110011000000011011;
#10000;
	data_in <= 24'b010100000011000100011100;
#10000;
	data_in <= 24'b010100110011001000011111;
#10000;
	data_in <= 24'b010101000011001000100010;
#10000;
	data_in <= 24'b010100110011001000100011;
#10000;
	data_in <= 24'b010011110011001000100100;
#10000;
	data_in <= 24'b010011100011010000100110;
#10000;
	data_in <= 24'b010100010011011100101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100100011100101010011;
#10000;
	data_in <= 24'b010000110011010001010100;
#10000;
	data_in <= 24'b010000010011101001011111;
#10000;
	data_in <= 24'b011000010101111110000011;
#10000;
	data_in <= 24'b100010001000010110100101;
#10000;
	data_in <= 24'b011010110110010001111111;
#10000;
	data_in <= 24'b010011010100000101010101;
#10000;
	data_in <= 24'b010010100011100001000101;
#10000;
	data_in <= 24'b010011010011010001001110;
#10000;
	data_in <= 24'b010010010011100001011010;
#10000;
	data_in <= 24'b010001100011111001100111;
#10000;
	data_in <= 24'b010100010100110101110110;
#10000;
	data_in <= 24'b100010011000010110101000;
#10000;
	data_in <= 24'b011010000110001110000000;
#10000;
	data_in <= 24'b010011010100000101010111;
#10000;
	data_in <= 24'b010001000011001101000001;
#10000;
	data_in <= 24'b010100000011100101001111;
#10000;
	data_in <= 24'b010100100011111101100000;
#10000;
	data_in <= 24'b010010100011110001100101;
#10000;
	data_in <= 24'b010011110100011001101110;
#10000;
	data_in <= 24'b010110100101001101110110;
#10000;
	data_in <= 24'b010110000101000001101110;
#10000;
	data_in <= 24'b010011100100000101011001;
#10000;
	data_in <= 24'b010010010011011101001000;
#10000;
	data_in <= 24'b010010010011001001000001;
#10000;
	data_in <= 24'b010011010011100001010001;
#10000;
	data_in <= 24'b010110000100011101101000;
#10000;
	data_in <= 24'b010101010100010101100111;
#10000;
	data_in <= 24'b010101010100011001100110;
#10000;
	data_in <= 24'b010010100011110001011000;
#10000;
	data_in <= 24'b010100000100001101011001;
#10000;
	data_in <= 24'b010001100011010001000101;
#10000;
	data_in <= 24'b010001110011000000110101;
#10000;
	data_in <= 24'b010011100011011101000101;
#10000;
	data_in <= 24'b010101010011111001010100;
#10000;
	data_in <= 24'b010110100100001001011010;
#10000;
	data_in <= 24'b011001100101000001101000;
#10000;
	data_in <= 24'b010110010100010001011010;
#10000;
	data_in <= 24'b010100110100000001010011;
#10000;
	data_in <= 24'b010011110011101001001001;
#10000;
	data_in <= 24'b010100010011101000111000;
#10000;
	data_in <= 24'b010100000011011100111011;
#10000;
	data_in <= 24'b010011010011000000111001;
#10000;
	data_in <= 24'b010111010011111101001100;
#10000;
	data_in <= 24'b010111010011111001001101;
#10000;
	data_in <= 24'b010111100100001101010011;
#10000;
	data_in <= 24'b010101100011111101001110;
#10000;
	data_in <= 24'b010101010011111001001101;
#10000;
	data_in <= 24'b010101000011101100110001;
#10000;
	data_in <= 24'b010011100011001000101011;
#10000;
	data_in <= 24'b010110100011100100110110;
#10000;
	data_in <= 24'b010110110011011000111000;
#10000;
	data_in <= 24'b010110110011010000111100;
#10000;
	data_in <= 24'b010100100010111000111010;
#10000;
	data_in <= 24'b010101110011101001001001;
#10000;
	data_in <= 24'b010010000010111000111100;
#10000;
	data_in <= 24'b010100100011100000101010;
#10000;
	data_in <= 24'b010111100100000100110011;
#10000;
	data_in <= 24'b010110000011010100101011;
#10000;
	data_in <= 24'b010101110011000100101100;
#10000;
	data_in <= 24'b010101100010111100101101;
#10000;
	data_in <= 24'b010101110011001000110100;
#10000;
	data_in <= 24'b010011110010111100110100;
#10000;
	data_in <= 24'b010010110010110100110010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010000100010101100110000;
#10000;
	data_in <= 24'b010001000010100100101100;
#10000;
	data_in <= 24'b010000110010011100100111;
#10000;
	data_in <= 24'b010001110010101100101010;
#10000;
	data_in <= 24'b010001100010101100100111;
#10000;
	data_in <= 24'b010000010010011100100001;
#10000;
	data_in <= 24'b010001000010100000100001;
#10000;
	data_in <= 24'b010001000010100000100001;
#10000;
	data_in <= 24'b010000110010101100110011;
#10000;
	data_in <= 24'b010001100010101100101111;
#10000;
	data_in <= 24'b010010000010101100101110;
#10000;
	data_in <= 24'b010010110010111100101111;
#10000;
	data_in <= 24'b010010010010110100101100;
#10000;
	data_in <= 24'b010001000010100100100101;
#10000;
	data_in <= 24'b010001010010100000100011;
#10000;
	data_in <= 24'b010001010010100100100010;
#10000;
	data_in <= 24'b010010000010111100111001;
#10000;
	data_in <= 24'b010010100010111000110100;
#10000;
	data_in <= 24'b010011000010111000110011;
#10000;
	data_in <= 24'b010011000010111100110010;
#10000;
	data_in <= 24'b010011000010110100101110;
#10000;
	data_in <= 24'b010010000010101000101001;
#10000;
	data_in <= 24'b010001110010100100100100;
#10000;
	data_in <= 24'b010001110010101000100011;
#10000;
	data_in <= 24'b010011010011001101000000;
#10000;
	data_in <= 24'b010011010011000000111001;
#10000;
	data_in <= 24'b010011100010111100110110;
#10000;
	data_in <= 24'b010010110010110100110010;
#10000;
	data_in <= 24'b010010110010110000101101;
#10000;
	data_in <= 24'b010010100010110000101011;
#10000;
	data_in <= 24'b010001100010100000100011;
#10000;
	data_in <= 24'b010001100010100100100010;
#10000;
	data_in <= 24'b010100010011011101000100;
#10000;
	data_in <= 24'b010100000011001100111100;
#10000;
	data_in <= 24'b010100100011001100111010;
#10000;
	data_in <= 24'b010011100011000000110101;
#10000;
	data_in <= 24'b010011110011000000110001;
#10000;
	data_in <= 24'b010100000011001100101111;
#10000;
	data_in <= 24'b010010000010101100100100;
#10000;
	data_in <= 24'b010001010010100000011111;
#10000;
	data_in <= 24'b010101010011100101000110;
#10000;
	data_in <= 24'b010100110011011000111111;
#10000;
	data_in <= 24'b010110010011101001000001;
#10000;
	data_in <= 24'b010101000011011000111011;
#10000;
	data_in <= 24'b010101100011011100111000;
#10000;
	data_in <= 24'b010110000011101100110111;
#10000;
	data_in <= 24'b010010110010111000100111;
#10000;
	data_in <= 24'b010001110010101100100000;
#10000;
	data_in <= 24'b010100000011010100111111;
#10000;
	data_in <= 24'b010011110011001000111011;
#10000;
	data_in <= 24'b010101110011100000111111;
#10000;
	data_in <= 24'b010100010011010000110111;
#10000;
	data_in <= 24'b010100100011010000110011;
#10000;
	data_in <= 24'b010101100011100100110100;
#10000;
	data_in <= 24'b010010100010110100100100;
#10000;
	data_in <= 24'b010010000010110000100001;
#10000;
	data_in <= 24'b010010100010110100110000;
#10000;
	data_in <= 24'b010010100010101100101100;
#10000;
	data_in <= 24'b010100010011001100110010;
#10000;
	data_in <= 24'b010010000010101100100111;
#10000;
	data_in <= 24'b010001110010101000100011;
#10000;
	data_in <= 24'b010011010011000000100111;
#10000;
	data_in <= 24'b010001100010100100011011;
#10000;
	data_in <= 24'b010010000010101100011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010000100010010100011100;
#10000;
	data_in <= 24'b010000100010010100011100;
#10000;
	data_in <= 24'b010000100010010100011100;
#10000;
	data_in <= 24'b010000010010010000011011;
#10000;
	data_in <= 24'b010000000010001100011010;
#10000;
	data_in <= 24'b001111100010000100011000;
#10000;
	data_in <= 24'b001110110001111000010111;
#10000;
	data_in <= 24'b001110000001110000010101;
#10000;
	data_in <= 24'b010000010010010000011011;
#10000;
	data_in <= 24'b010000010010010000011011;
#10000;
	data_in <= 24'b010000010010010000011011;
#10000;
	data_in <= 24'b010000010010010000011011;
#10000;
	data_in <= 24'b010000000010001100011010;
#10000;
	data_in <= 24'b001111100010000100011000;
#10000;
	data_in <= 24'b001110110001111000010111;
#10000;
	data_in <= 24'b001110100001110100010110;
#10000;
	data_in <= 24'b010000010010001000011001;
#10000;
	data_in <= 24'b010000100010001100011010;
#10000;
	data_in <= 24'b010000100010010000011001;
#10000;
	data_in <= 24'b010000100010010000011001;
#10000;
	data_in <= 24'b010000010010001100011000;
#10000;
	data_in <= 24'b001111110010000100010110;
#10000;
	data_in <= 24'b001111010001111000010101;
#10000;
	data_in <= 24'b001111000001110100010100;
#10000;
	data_in <= 24'b010000100010001100011010;
#10000;
	data_in <= 24'b010000110010010100011010;
#10000;
	data_in <= 24'b010000110010010100011010;
#10000;
	data_in <= 24'b010000100010010100010111;
#10000;
	data_in <= 24'b010000000010001100010101;
#10000;
	data_in <= 24'b001111100010000100010011;
#10000;
	data_in <= 24'b001111010001111100010100;
#10000;
	data_in <= 24'b001111010001111100010100;
#10000;
	data_in <= 24'b010001000010011000011011;
#10000;
	data_in <= 24'b010001000010011100011001;
#10000;
	data_in <= 24'b010001000010011100011001;
#10000;
	data_in <= 24'b010000110010011000010111;
#10000;
	data_in <= 24'b010000110010010000010101;
#10000;
	data_in <= 24'b010000010010001000010011;
#10000;
	data_in <= 24'b010000000010000000010011;
#10000;
	data_in <= 24'b001111110001111100010010;
#10000;
	data_in <= 24'b010001110010101000011100;
#10000;
	data_in <= 24'b010001010010100000011001;
#10000;
	data_in <= 24'b010001000010011100011000;
#10000;
	data_in <= 24'b010000110010011100010110;
#10000;
	data_in <= 24'b010001000010011000010101;
#10000;
	data_in <= 24'b010000100010010000010011;
#10000;
	data_in <= 24'b010000010010001100010010;
#10000;
	data_in <= 24'b001111110010000100010000;
#10000;
	data_in <= 24'b010010000010101100011100;
#10000;
	data_in <= 24'b010001010010100100011000;
#10000;
	data_in <= 24'b010001010010011100010100;
#10000;
	data_in <= 24'b010001000010011000010011;
#10000;
	data_in <= 24'b010001010010011100010100;
#10000;
	data_in <= 24'b010001000010011000010011;
#10000;
	data_in <= 24'b010000100010010000010001;
#10000;
	data_in <= 24'b010000000010001000001111;
#10000;
	data_in <= 24'b010010000010110000011011;
#10000;
	data_in <= 24'b010001110010100100010110;
#10000;
	data_in <= 24'b010001000010011100010010;
#10000;
	data_in <= 24'b010001000010011100010010;
#10000;
	data_in <= 24'b010001010010100000010011;
#10000;
	data_in <= 24'b010001010010100000010011;
#10000;
	data_in <= 24'b010000110010011000010001;
#10000;
	data_in <= 24'b010000000010001100001110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001000110001000000001011;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b001010000001010100010000;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001011000001100100010010;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001000010000111000001001;
#10000;
	data_in <= 24'b001000110001000000001011;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001001110001010000001111;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001011000001100100010010;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001000100000111100001010;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b001010000001010100010000;
#10000;
	data_in <= 24'b001010110001100100010010;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001000110001000000001011;
#10000;
	data_in <= 24'b001001110001010000001111;
#10000;
	data_in <= 24'b001010000001010100010000;
#10000;
	data_in <= 24'b001010010001011000010001;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b001011010001101100010100;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001001000001000100001100;
#10000;
	data_in <= 24'b001001110001010000001111;
#10000;
	data_in <= 24'b001010000001010100010000;
#10000;
	data_in <= 24'b001010010001011000010001;
#10000;
	data_in <= 24'b001010110001100100010010;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001010010001011000010001;
#10000;
	data_in <= 24'b001010100001011100010010;
#10000;
	data_in <= 24'b001010100001011100010010;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b001011010001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b001010110001100000010011;
#10000;
	data_in <= 24'b001010110001100100010010;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001001010001001000001101;
#10000;
	data_in <= 24'b001010010001011000010001;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001010010001011100010000;
#10000;
	data_in <= 24'b001011010001101000010011;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001101010010001000011011;
#10000;
	data_in <= 24'b001110000010010100011101;
#10000;
	data_in <= 24'b001110100010011100011111;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001101100010001100011100;
#10000;
	data_in <= 24'b001110010010011000011110;
#10000;
	data_in <= 24'b001110100010011100011111;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001101100010001100011100;
#10000;
	data_in <= 24'b001110010010011000011110;
#10000;
	data_in <= 24'b001110110010100000100000;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000010010110000100100;
#10000;
	data_in <= 24'b010000010010110000100100;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001101100010001100011100;
#10000;
	data_in <= 24'b001110000010010100011101;
#10000;
	data_in <= 24'b001110100010011100011111;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b010000010010110000100100;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b001100110010000000011000;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001101100010001100011011;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001101110010010000011100;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b001111010010100100011110;
#10000;
	data_in <= 24'b001101110010010000011100;
#10000;
	data_in <= 24'b001110000010010100011101;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b001111010010100100011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010000000010100100100001;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000000010101000011110;
#10000;
	data_in <= 24'b010000100010110000100000;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b010001010011000000100001;
#10000;
	data_in <= 24'b010000110010111000011111;
#10000;
	data_in <= 24'b010000110010110000100100;
#10000;
	data_in <= 24'b010000110010110000100100;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010001010010111100100011;
#10000;
	data_in <= 24'b010010000011001000100110;
#10000;
	data_in <= 24'b010010010011010000100101;
#10000;
	data_in <= 24'b010010000011001100100100;
#10000;
	data_in <= 24'b010000110010110000100100;
#10000;
	data_in <= 24'b010001000010110100100101;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001100011000000100100;
#10000;
	data_in <= 24'b010010010011001100100111;
#10000;
	data_in <= 24'b010011010011011000100111;
#10000;
	data_in <= 24'b010011100011011100101000;
#10000;
	data_in <= 24'b010000100010101100100011;
#10000;
	data_in <= 24'b010000110010110000100100;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b010001100011000000100100;
#10000;
	data_in <= 24'b010010110011010000100101;
#10000;
	data_in <= 24'b010011010011011000100111;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010000110010110100100001;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b010010010011001000100011;
#10000;
	data_in <= 24'b010010110011010000100101;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000110010110100100001;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b010010000011000100100010;
#10000;
	data_in <= 24'b010010100011001100100100;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010001010010110100100001;
#10000;
	data_in <= 24'b010001110010111100100011;
#10000;
	data_in <= 24'b010001110011000000100001;
#10000;
	data_in <= 24'b010001110011000000100001;
#10000;
	data_in <= 24'b010010010011001000100011;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b001111100010100000011101;
#10000;
	data_in <= 24'b010000010010100100011101;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010001110011000000100001;
#10000;
	data_in <= 24'b010001110011000000100001;
#10000;
	data_in <= 24'b010001100010111100100000;
#10000;
	data_in <= 24'b010001110011000000100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010010010011001000100011;
#10000;
	data_in <= 24'b010010110011010000100101;
#10000;
	data_in <= 24'b010011010011011000100110;
#10000;
	data_in <= 24'b010011110011100000101000;
#10000;
	data_in <= 24'b010011100011011100100111;
#10000;
	data_in <= 24'b010011100011011100100111;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010011000011010100100110;
#10000;
	data_in <= 24'b010011100011011100101000;
#10000;
	data_in <= 24'b010100000011100100101001;
#10000;
	data_in <= 24'b010100100011101100101011;
#10000;
	data_in <= 24'b010100100011101100101011;
#10000;
	data_in <= 24'b010100010011101000101010;
#10000;
	data_in <= 24'b010100010011100000101000;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010100000011100100101001;
#10000;
	data_in <= 24'b010100010011101000101010;
#10000;
	data_in <= 24'b010100110011110000101100;
#10000;
	data_in <= 24'b010101010011111000101110;
#10000;
	data_in <= 24'b010101110011111000101110;
#10000;
	data_in <= 24'b010101100011110100101101;
#10000;
	data_in <= 24'b010100110011101000101010;
#10000;
	data_in <= 24'b010100010011100000101000;
#10000;
	data_in <= 24'b010100100011101100101011;
#10000;
	data_in <= 24'b010100100011101100101011;
#10000;
	data_in <= 24'b010100110011110000101100;
#10000;
	data_in <= 24'b010101000011110100101101;
#10000;
	data_in <= 24'b010101110011111000101110;
#10000;
	data_in <= 24'b010101110011111000101110;
#10000;
	data_in <= 24'b010101000011101100101011;
#10000;
	data_in <= 24'b010100100011100100101001;
#10000;
	data_in <= 24'b010100000011100100101001;
#10000;
	data_in <= 24'b010100000011100100101001;
#10000;
	data_in <= 24'b010100100011100100101001;
#10000;
	data_in <= 24'b010100110011101000101010;
#10000;
	data_in <= 24'b010101010011110000101100;
#10000;
	data_in <= 24'b010101010011110000101100;
#10000;
	data_in <= 24'b010101000011101000101100;
#10000;
	data_in <= 24'b010100110011101000101010;
#10000;
	data_in <= 24'b010011010011011000100110;
#10000;
	data_in <= 24'b010011010011011000100110;
#10000;
	data_in <= 24'b010011110011011000100110;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010100010011100000101000;
#10000;
	data_in <= 24'b010100110011101000101010;
#10000;
	data_in <= 24'b010100110011100100101011;
#10000;
	data_in <= 24'b010100110011100100101011;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010011010011010000100100;
#10000;
	data_in <= 24'b010011100011010100100101;
#10000;
	data_in <= 24'b010011110011011000100110;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010100010011100000101000;
#10000;
	data_in <= 24'b010100010011011100101001;
#10000;
	data_in <= 24'b010100100011100000101010;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010011110011011000100110;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010100000011011100100111;
#10000;
	data_in <= 24'b010100000011011000101000;
#10000;
	data_in <= 24'b010100010011011100101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100100011100000101000;
#10000;
	data_in <= 24'b010011100011010000100011;
#10000;
	data_in <= 24'b010011100011010000100011;
#10000;
	data_in <= 24'b010011000011001000100001;
#10000;
	data_in <= 24'b010010010010111100011110;
#10000;
	data_in <= 24'b010011010011001100100010;
#10000;
	data_in <= 24'b010100000011010000100011;
#10000;
	data_in <= 24'b010010010010110100011100;
#10000;
	data_in <= 24'b010100010011011100100110;
#10000;
	data_in <= 24'b010011010011001100100010;
#10000;
	data_in <= 24'b010011010011001100100010;
#10000;
	data_in <= 24'b010010110011000100100000;
#10000;
	data_in <= 24'b010010000010111000011101;
#10000;
	data_in <= 24'b010010100011000000011111;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010011000011000000011111;
#10000;
	data_in <= 24'b010100010011011100100110;
#10000;
	data_in <= 24'b010011010011001100100010;
#10000;
	data_in <= 24'b010011000011001000100001;
#10000;
	data_in <= 24'b010010110011000100100000;
#10000;
	data_in <= 24'b010001110010110100011100;
#10000;
	data_in <= 24'b010001110010110100011100;
#10000;
	data_in <= 24'b010011010011000100100000;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010100100011100000101000;
#10000;
	data_in <= 24'b010011100011010000100011;
#10000;
	data_in <= 24'b010010110011000100100000;
#10000;
	data_in <= 24'b010010110011000100100000;
#10000;
	data_in <= 24'b010010010010111100011110;
#10000;
	data_in <= 24'b010001110010110100011100;
#10000;
	data_in <= 24'b010010110010111100011110;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010101000011101000101010;
#10000;
	data_in <= 24'b010011110011010100100101;
#10000;
	data_in <= 24'b010011000011001000100001;
#10000;
	data_in <= 24'b010011010011001100100010;
#10000;
	data_in <= 24'b010011010011001100100010;
#10000;
	data_in <= 24'b010010000010111000011101;
#10000;
	data_in <= 24'b010010010010111000011010;
#10000;
	data_in <= 24'b010011010011001000011110;
#10000;
	data_in <= 24'b010101000011101000101010;
#10000;
	data_in <= 24'b010100010011011100100111;
#10000;
	data_in <= 24'b010011100011010000100011;
#10000;
	data_in <= 24'b010011100011010000100011;
#10000;
	data_in <= 24'b010100000011011000100101;
#10000;
	data_in <= 24'b010010110011000100100000;
#10000;
	data_in <= 24'b010010100010111100011011;
#10000;
	data_in <= 24'b010011010011001000011110;
#10000;
	data_in <= 24'b010100100011100000101000;
#10000;
	data_in <= 24'b010101000011101000101010;
#10000;
	data_in <= 24'b010100010011011100100111;
#10000;
	data_in <= 24'b010100000011011000100110;
#10000;
	data_in <= 24'b010100110011011100100110;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010011000011000100011101;
#10000;
	data_in <= 24'b010100000011010100100001;
#10000;
	data_in <= 24'b010100010011011100100111;
#10000;
	data_in <= 24'b010101010011101100101011;
#10000;
	data_in <= 24'b010100110011100100101001;
#10000;
	data_in <= 24'b010100000011011000100110;
#10000;
	data_in <= 24'b010100110011011100100110;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010011100011001100011111;
#10000;
	data_in <= 24'b010101000011100100100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010011000011000000011111;
#10000;
	data_in <= 24'b010011000011000100011101;
#10000;
	data_in <= 24'b010010110010110100011100;
#10000;
	data_in <= 24'b010010110010110100011010;
#10000;
	data_in <= 24'b010011110011000100100000;
#10000;
	data_in <= 24'b010011110011000100011110;
#10000;
	data_in <= 24'b010010110010110100011100;
#10000;
	data_in <= 24'b010011000010110000011001;
#10000;
	data_in <= 24'b010010100010111000011101;
#10000;
	data_in <= 24'b010010110010111100011110;
#10000;
	data_in <= 24'b010010110010110100011100;
#10000;
	data_in <= 24'b010011000010111000011101;
#10000;
	data_in <= 24'b010011110011000100100000;
#10000;
	data_in <= 24'b010011110011000100100000;
#10000;
	data_in <= 24'b010011010010110000011100;
#10000;
	data_in <= 24'b010011000010110000011001;
#10000;
	data_in <= 24'b010010000010110100011001;
#10000;
	data_in <= 24'b010010100010111100011011;
#10000;
	data_in <= 24'b010011000010111000011011;
#10000;
	data_in <= 24'b010011010010111100011100;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100010011000100011110;
#10000;
	data_in <= 24'b010011100010111000011011;
#10000;
	data_in <= 24'b010011100010111000011011;
#10000;
	data_in <= 24'b010010010010111000011010;
#10000;
	data_in <= 24'b010010110011000000011100;
#10000;
	data_in <= 24'b010011010010111100011100;
#10000;
	data_in <= 24'b010011100011000000011101;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100000011000000011101;
#10000;
	data_in <= 24'b010011110010111100011100;
#10000;
	data_in <= 24'b010100010011001000011101;
#10000;
	data_in <= 24'b010011010010111100011100;
#10000;
	data_in <= 24'b010011100011000000011101;
#10000;
	data_in <= 24'b010011010011000000011011;
#10000;
	data_in <= 24'b010011100011000100011100;
#10000;
	data_in <= 24'b010100100011001100011110;
#10000;
	data_in <= 24'b010100000011000100011100;
#10000;
	data_in <= 24'b010100000011000100011100;
#10000;
	data_in <= 24'b010101000011010100100000;
#10000;
	data_in <= 24'b010100000011001000011111;
#10000;
	data_in <= 24'b010100000011001000011111;
#10000;
	data_in <= 24'b010011100011000100011100;
#10000;
	data_in <= 24'b010011110011001000011101;
#10000;
	data_in <= 24'b010100110011010000011111;
#10000;
	data_in <= 24'b010100010011001000011101;
#10000;
	data_in <= 24'b010100010011001000011101;
#10000;
	data_in <= 24'b010101010011011000100001;
#10000;
	data_in <= 24'b010100110011010100100010;
#10000;
	data_in <= 24'b010100010011001100100000;
#10000;
	data_in <= 24'b010011110011001000011101;
#10000;
	data_in <= 24'b010100010011010000011111;
#10000;
	data_in <= 24'b010101010011011000011111;
#10000;
	data_in <= 24'b010100100011001100011100;
#10000;
	data_in <= 24'b010100010011001000011011;
#10000;
	data_in <= 24'b010101010011011000011111;
#10000;
	data_in <= 24'b010101000011011000100011;
#10000;
	data_in <= 24'b010100100011010000100001;
#10000;
	data_in <= 24'b010100000011001100011110;
#10000;
	data_in <= 24'b010100100011010100100000;
#10000;
	data_in <= 24'b010101110011100000100001;
#10000;
	data_in <= 24'b010101000011010100011110;
#10000;
	data_in <= 24'b010100010011001000011011;
#10000;
	data_in <= 24'b010101000011010100011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010010100010101100010110;
#10000;
	data_in <= 24'b010010110010110000010111;
#10000;
	data_in <= 24'b010010110010110000010111;
#10000;
	data_in <= 24'b010010100010100100010101;
#10000;
	data_in <= 24'b010011010010110000011000;
#10000;
	data_in <= 24'b010101000011000100011101;
#10000;
	data_in <= 24'b010100110010111100011101;
#10000;
	data_in <= 24'b010011110010101100011001;
#10000;
	data_in <= 24'b010010110010110000010111;
#10000;
	data_in <= 24'b010100000011000100011100;
#10000;
	data_in <= 24'b010100000011000100011100;
#10000;
	data_in <= 24'b010011000010110100011000;
#10000;
	data_in <= 24'b010011100010110100011001;
#10000;
	data_in <= 24'b010100100011000100011101;
#10000;
	data_in <= 24'b010101000011000000011110;
#10000;
	data_in <= 24'b010011110010101100011001;
#10000;
	data_in <= 24'b010011010010111000011001;
#10000;
	data_in <= 24'b010100110011010000011101;
#10000;
	data_in <= 24'b010101000011001100011111;
#10000;
	data_in <= 24'b010011110010111000011010;
#10000;
	data_in <= 24'b010011100010110100011001;
#10000;
	data_in <= 24'b010100110011001000011110;
#10000;
	data_in <= 24'b010101010011001000011110;
#10000;
	data_in <= 24'b010100010010111000011010;
#10000;
	data_in <= 24'b010100000011000100011010;
#10000;
	data_in <= 24'b010100010011001000011011;
#10000;
	data_in <= 24'b010100100011000100011101;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010100100011000100011101;
#10000;
	data_in <= 24'b010101010011001000011110;
#10000;
	data_in <= 24'b010101000011000100011101;
#10000;
	data_in <= 24'b010101100011011000011111;
#10000;
	data_in <= 24'b010100100011001000011011;
#10000;
	data_in <= 24'b010011110010111100011000;
#10000;
	data_in <= 24'b010100000011000000011001;
#10000;
	data_in <= 24'b010101000011001000011011;
#10000;
	data_in <= 24'b010100110011000100011010;
#10000;
	data_in <= 24'b010100110011000000011100;
#10000;
	data_in <= 24'b010101010011001000011110;
#10000;
	data_in <= 24'b010110100011101000100011;
#10000;
	data_in <= 24'b010101000011010000011101;
#10000;
	data_in <= 24'b010100010011000100011010;
#10000;
	data_in <= 24'b010100110011001100011100;
#10000;
	data_in <= 24'b010101100011010000011101;
#10000;
	data_in <= 24'b010101000011001000011011;
#10000;
	data_in <= 24'b010100110011000000011100;
#10000;
	data_in <= 24'b010100110011000000011100;
#10000;
	data_in <= 24'b010101110011011100100000;
#10000;
	data_in <= 24'b010101110011011100100000;
#10000;
	data_in <= 24'b010101100011011000011111;
#10000;
	data_in <= 24'b010101010011010100011110;
#10000;
	data_in <= 24'b010101100011010000011101;
#10000;
	data_in <= 24'b010101100011010000011101;
#10000;
	data_in <= 24'b010101000011001000011011;
#10000;
	data_in <= 24'b010100010010111100011000;
#10000;
	data_in <= 24'b010100100011001000011011;
#10000;
	data_in <= 24'b010110000011100000100001;
#10000;
	data_in <= 24'b010110100011101000100011;
#10000;
	data_in <= 24'b010101010011010100011110;
#10000;
	data_in <= 24'b010101100011010000011101;
#10000;
	data_in <= 24'b010110000011011000011111;
#10000;
	data_in <= 24'b010101100011010000011101;
#10000;
	data_in <= 24'b010100000010111000010111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100110010111100011101;
#10000;
	data_in <= 24'b010101000011000000011110;
#10000;
	data_in <= 24'b010100110010111100011101;
#10000;
	data_in <= 24'b010100010010110100011011;
#10000;
	data_in <= 24'b010100100010111000011100;
#10000;
	data_in <= 24'b010101100011001100011111;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010100100011000100011101;
#10000;
	data_in <= 24'b010101100011001000100000;
#10000;
	data_in <= 24'b010101010011000100011111;
#10000;
	data_in <= 24'b010101000011000000011110;
#10000;
	data_in <= 24'b010100110010111100011101;
#10000;
	data_in <= 24'b010100110010111100011101;
#10000;
	data_in <= 24'b010101010011000100011111;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010100110011001000011111;
#10000;
	data_in <= 24'b010101100011001000100000;
#10000;
	data_in <= 24'b010101100011001000100000;
#10000;
	data_in <= 24'b010101110011001100100001;
#10000;
	data_in <= 24'b010110010011010100100011;
#10000;
	data_in <= 24'b010101100011010100100010;
#10000;
	data_in <= 24'b010101010011010000100001;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010101010011010000100001;
#10000;
	data_in <= 24'b010101000011000000011110;
#10000;
	data_in <= 24'b010101100011001000100000;
#10000;
	data_in <= 24'b010110100011011000100100;
#10000;
	data_in <= 24'b010111100011101000101000;
#10000;
	data_in <= 24'b010110110011101000100111;
#10000;
	data_in <= 24'b010101110011011000100011;
#10000;
	data_in <= 24'b010101010011010000100001;
#10000;
	data_in <= 24'b010101100011010100100010;
#10000;
	data_in <= 24'b010101000011000100011101;
#10000;
	data_in <= 24'b010101100011001100011111;
#10000;
	data_in <= 24'b010110000011011100100100;
#10000;
	data_in <= 24'b010110110011101000100111;
#10000;
	data_in <= 24'b010110110011101000100111;
#10000;
	data_in <= 24'b010101100011010100100010;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100110011001100100000;
#10000;
	data_in <= 24'b010101100011001100011111;
#10000;
	data_in <= 24'b010101110011010000100000;
#10000;
	data_in <= 24'b010101110011011000100011;
#10000;
	data_in <= 24'b010110000011011100100100;
#10000;
	data_in <= 24'b010101110011011000100011;
#10000;
	data_in <= 24'b010101010011010000100001;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010101110011010000100000;
#10000;
	data_in <= 24'b010110100011011100100011;
#10000;
	data_in <= 24'b010110100011100100100101;
#10000;
	data_in <= 24'b010110110011101000100110;
#10000;
	data_in <= 24'b010110110011101000100111;
#10000;
	data_in <= 24'b010110100011100100100110;
#10000;
	data_in <= 24'b010101100011010100100101;
#10000;
	data_in <= 24'b010100110011001000100010;
#10000;
	data_in <= 24'b010101100011001100011111;
#10000;
	data_in <= 24'b010110110011100000100100;
#10000;
	data_in <= 24'b010111100011110100101001;
#10000;
	data_in <= 24'b011000010100000000101100;
#10000;
	data_in <= 24'b011000110100001000101111;
#10000;
	data_in <= 24'b011000100100000100101110;
#10000;
	data_in <= 24'b010111000011101100101011;
#10000;
	data_in <= 24'b010101100011010100100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010011110010111100011100;
#10000;
	data_in <= 24'b010100010011000100011110;
#10000;
	data_in <= 24'b010101000011010000100001;
#10000;
	data_in <= 24'b010101110011011000100110;
#10000;
	data_in <= 24'b010101000011011000100101;
#10000;
	data_in <= 24'b010100110011010000100101;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100110011001100100000;
#10000;
	data_in <= 24'b010100110011001100100000;
#10000;
	data_in <= 24'b010100110011010100100010;
#10000;
	data_in <= 24'b010101000011011000100011;
#10000;
	data_in <= 24'b010100110011010100100100;
#10000;
	data_in <= 24'b010100010011001100100010;
#10000;
	data_in <= 24'b010100000011001000100001;
#10000;
	data_in <= 24'b010100100011010000100011;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100110011001100100000;
#10000;
	data_in <= 24'b010101000011010000100001;
#10000;
	data_in <= 24'b010101010011010100100010;
#10000;
	data_in <= 24'b010101000011001100100011;
#10000;
	data_in <= 24'b010100100011000100100001;
#10000;
	data_in <= 24'b010100110011001000100010;
#10000;
	data_in <= 24'b010101000011001100100011;
#10000;
	data_in <= 24'b010100010011000100011110;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100110011001100100000;
#10000;
	data_in <= 24'b010101000011010000100001;
#10000;
	data_in <= 24'b010101000011001100100011;
#10000;
	data_in <= 24'b010100100011000100100001;
#10000;
	data_in <= 24'b010100110011001000100010;
#10000;
	data_in <= 24'b010101000011010000100001;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010100110011001000011111;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010101010011010000100001;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010100010011000000011101;
#10000;
	data_in <= 24'b010100010011000000011101;
#10000;
	data_in <= 24'b010100010011000000011101;
#10000;
	data_in <= 24'b010100110011001000011111;
#10000;
	data_in <= 24'b010100110011001000011111;
#10000;
	data_in <= 24'b010100110011001000011111;
#10000;
	data_in <= 24'b010101010011010000100001;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010100100011000100011110;
#10000;
	data_in <= 24'b010100010011000000011101;
#10000;
	data_in <= 24'b010100110011000000011100;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010101110011001100100001;
#10000;
	data_in <= 24'b010110010011010100100011;
#10000;
	data_in <= 24'b010110010011010100100011;
#10000;
	data_in <= 24'b010101110011001100100001;
#10000;
	data_in <= 24'b010101010011001000011110;
#10000;
	data_in <= 24'b010101010011001000011110;
#10000;
	data_in <= 24'b010110100011100100100110;
#10000;
	data_in <= 24'b010110010011100000100101;
#10000;
	data_in <= 24'b010111000011100000100110;
#10000;
	data_in <= 24'b010111010011100100100111;
#10000;
	data_in <= 24'b010111000011100000100110;
#10000;
	data_in <= 24'b010110010011010100100011;
#10000;
	data_in <= 24'b010101010011001000011110;
#10000;
	data_in <= 24'b010101100011000100011101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010101110011100100101000;
#10000;
	data_in <= 24'b010101110011100000101001;
#10000;
	data_in <= 24'b010101110011011000100111;
#10000;
	data_in <= 24'b010101010011001100100110;
#10000;
	data_in <= 24'b010101000011001000100101;
#10000;
	data_in <= 24'b010100000011000000100011;
#10000;
	data_in <= 24'b010011000010111100100001;
#10000;
	data_in <= 24'b010101000011011000100101;
#10000;
	data_in <= 24'b010101000011011000100011;
#10000;
	data_in <= 24'b010101000011011000100011;
#10000;
	data_in <= 24'b010100110011001100100000;
#10000;
	data_in <= 24'b010100010011000100011110;
#10000;
	data_in <= 24'b010100000011000100011100;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010011100010110100011001;
#10000;
	data_in <= 24'b010101000011010000100001;
#10000;
	data_in <= 24'b010101000011010000100001;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100000010111100011011;
#10000;
	data_in <= 24'b010011110010111000011010;
#10000;
	data_in <= 24'b010011100010110100011001;
#10000;
	data_in <= 24'b010011110010110000011000;
#10000;
	data_in <= 24'b010011100010110000010101;
#10000;
	data_in <= 24'b010101010011010100100010;
#10000;
	data_in <= 24'b010101000011001100011111;
#10000;
	data_in <= 24'b010100100011000100011101;
#10000;
	data_in <= 24'b010100010010111000011010;
#10000;
	data_in <= 24'b010100000010110100011001;
#10000;
	data_in <= 24'b010100100010110100010111;
#10000;
	data_in <= 24'b010100100010110100010111;
#10000;
	data_in <= 24'b010100010010110100010101;
#10000;
	data_in <= 24'b010101000011001100100000;
#10000;
	data_in <= 24'b010101000011000100011101;
#10000;
	data_in <= 24'b010100100010111100011011;
#10000;
	data_in <= 24'b010100110010111000011000;
#10000;
	data_in <= 24'b010100110010111000011000;
#10000;
	data_in <= 24'b010101010010111100010111;
#10000;
	data_in <= 24'b010101000010111000010110;
#10000;
	data_in <= 24'b010101000010111100010101;
#10000;
	data_in <= 24'b010101010011001000011110;
#10000;
	data_in <= 24'b010101000010111100011001;
#10000;
	data_in <= 24'b010100110010111000011000;
#10000;
	data_in <= 24'b010101010010111100010111;
#10000;
	data_in <= 24'b010101010010111100010111;
#10000;
	data_in <= 24'b010101110010111100010110;
#10000;
	data_in <= 24'b010101100010111000010101;
#10000;
	data_in <= 24'b010101110010111000010101;
#10000;
	data_in <= 24'b010101110011001000011110;
#10000;
	data_in <= 24'b010101110011000000011010;
#10000;
	data_in <= 24'b010101100011000000011000;
#10000;
	data_in <= 24'b010110010011000100011000;
#10000;
	data_in <= 24'b010110100011001000011001;
#10000;
	data_in <= 24'b010110010011000100010101;
#10000;
	data_in <= 24'b010101110010111100010011;
#10000;
	data_in <= 24'b010110010010111000010011;
#10000;
	data_in <= 24'b010110110011010000011110;
#10000;
	data_in <= 24'b010110010011001100011011;
#10000;
	data_in <= 24'b010110110011001100011010;
#10000;
	data_in <= 24'b010111000011010100011001;
#10000;
	data_in <= 24'b010111100011011000011010;
#10000;
	data_in <= 24'b010110110011001100010110;
#10000;
	data_in <= 24'b010110110011000100010100;
#10000;
	data_in <= 24'b010110100011000000010011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010010010010110000011101;
#10000;
	data_in <= 24'b010011010010111000011111;
#10000;
	data_in <= 24'b010011100010111100100000;
#10000;
	data_in <= 24'b010011110011000100100000;
#10000;
	data_in <= 24'b010100010011000000100000;
#10000;
	data_in <= 24'b010011110010111100011100;
#10000;
	data_in <= 24'b010010110010101100011000;
#10000;
	data_in <= 24'b010001110010100000010011;
#10000;
	data_in <= 24'b010011100010111000010111;
#10000;
	data_in <= 24'b010100010011000100011010;
#10000;
	data_in <= 24'b010100100011001000011011;
#10000;
	data_in <= 24'b010100010011000100011010;
#10000;
	data_in <= 24'b010011110010111100011000;
#10000;
	data_in <= 24'b010011010010110100010110;
#10000;
	data_in <= 24'b010011100010110000010101;
#10000;
	data_in <= 24'b010010100010101000010011;
#10000;
	data_in <= 24'b010011110010110100010110;
#10000;
	data_in <= 24'b010100110011000100011010;
#10000;
	data_in <= 24'b010101000011001000011010;
#10000;
	data_in <= 24'b010100010010111100010111;
#10000;
	data_in <= 24'b010011010010101100010011;
#10000;
	data_in <= 24'b010011000010101000010010;
#10000;
	data_in <= 24'b010011110010101100010011;
#10000;
	data_in <= 24'b010011100010110000010100;
#10000;
	data_in <= 24'b010100100010101100010101;
#10000;
	data_in <= 24'b010101010010111100010111;
#10000;
	data_in <= 24'b010101100011000000011000;
#10000;
	data_in <= 24'b010100110010110100010101;
#10000;
	data_in <= 24'b010100000010101000010010;
#10000;
	data_in <= 24'b010011110010100100010001;
#10000;
	data_in <= 24'b010100000010101000010010;
#10000;
	data_in <= 24'b010011110010101100010011;
#10000;
	data_in <= 24'b010100110010101000010011;
#10000;
	data_in <= 24'b010101010010110100010100;
#10000;
	data_in <= 24'b010101010010110100010100;
#10000;
	data_in <= 24'b010101000010110000010011;
#10000;
	data_in <= 24'b010100110010101100010010;
#10000;
	data_in <= 24'b010100110010101100010010;
#10000;
	data_in <= 24'b010100110010101100010010;
#10000;
	data_in <= 24'b010100000010101100010001;
#10000;
	data_in <= 24'b010101000010101100010010;
#10000;
	data_in <= 24'b010101010010110000010011;
#10000;
	data_in <= 24'b010101010010110000010011;
#10000;
	data_in <= 24'b010101010010110000010011;
#10000;
	data_in <= 24'b010101100010110100010100;
#10000;
	data_in <= 24'b010101100010110100010100;
#10000;
	data_in <= 24'b010101010010110000010011;
#10000;
	data_in <= 24'b010100010010100100010000;
#10000;
	data_in <= 24'b010110000010110100010010;
#10000;
	data_in <= 24'b010110010010111000010011;
#10000;
	data_in <= 24'b010110010010111000010011;
#10000;
	data_in <= 24'b010110000010110100010010;
#10000;
	data_in <= 24'b010110000010110100010010;
#10000;
	data_in <= 24'b010101110010111100010011;
#10000;
	data_in <= 24'b010101100010111000010010;
#10000;
	data_in <= 24'b010100110010101100001111;
#10000;
	data_in <= 24'b010110100010111100010100;
#10000;
	data_in <= 24'b010110110011000000010101;
#10000;
	data_in <= 24'b010110100010111100010100;
#10000;
	data_in <= 24'b010110010010111000010011;
#10000;
	data_in <= 24'b010110000010110100010010;
#10000;
	data_in <= 24'b010101110010111100010011;
#10000;
	data_in <= 24'b010101100010111000010010;
#10000;
	data_in <= 24'b010101000010110100010001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010001110010100000010011;
#10000;
	data_in <= 24'b010001010010011000010001;
#10000;
	data_in <= 24'b010001000010010100010000;
#10000;
	data_in <= 24'b010001000010010100010000;
#10000;
	data_in <= 24'b010000100010010000010001;
#10000;
	data_in <= 24'b010000010010001100010000;
#10000;
	data_in <= 24'b010000010010001100010000;
#10000;
	data_in <= 24'b010000110010010100010010;
#10000;
	data_in <= 24'b010010100010101000010011;
#10000;
	data_in <= 24'b010010000010100000010001;
#10000;
	data_in <= 24'b010001110010011000010010;
#10000;
	data_in <= 24'b010001100010011100010010;
#10000;
	data_in <= 24'b010001010010010100010010;
#10000;
	data_in <= 24'b010000010010001100010000;
#10000;
	data_in <= 24'b010000000010001000001111;
#10000;
	data_in <= 24'b010000000010001000001111;
#10000;
	data_in <= 24'b010010010010011100001111;
#10000;
	data_in <= 24'b010010010010011100001111;
#10000;
	data_in <= 24'b010010010010011100010000;
#10000;
	data_in <= 24'b010010000010100000010001;
#10000;
	data_in <= 24'b010010000010011100010011;
#10000;
	data_in <= 24'b010001010010011000010001;
#10000;
	data_in <= 24'b010000110010001100010000;
#10000;
	data_in <= 24'b010001000010010000010001;
#10000;
	data_in <= 24'b010011010010011100001111;
#10000;
	data_in <= 24'b010010110010011100001111;
#10000;
	data_in <= 24'b010010110010011000010000;
#10000;
	data_in <= 24'b010010100010100000010001;
#10000;
	data_in <= 24'b010010100010011100010011;
#10000;
	data_in <= 24'b010001110010011000010010;
#10000;
	data_in <= 24'b010001100010010100010010;
#10000;
	data_in <= 24'b010001100010011000010011;
#10000;
	data_in <= 24'b010100110010101100010010;
#10000;
	data_in <= 24'b010100000010101100010001;
#10000;
	data_in <= 24'b010011110010100100010001;
#10000;
	data_in <= 24'b010011010010100100010001;
#10000;
	data_in <= 24'b010010100010100000010001;
#10000;
	data_in <= 24'b010010000010011000001111;
#10000;
	data_in <= 24'b010001110010010000010000;
#10000;
	data_in <= 24'b010001100010010100010001;
#10000;
	data_in <= 24'b010101000010110000010011;
#10000;
	data_in <= 24'b010100100010101000010001;
#10000;
	data_in <= 24'b010100000010101000010010;
#10000;
	data_in <= 24'b010100000010101000010010;
#10000;
	data_in <= 24'b010011010010100000010010;
#10000;
	data_in <= 24'b010010100010100000010001;
#10000;
	data_in <= 24'b010010100010011100010011;
#10000;
	data_in <= 24'b010010110010100000010100;
#10000;
	data_in <= 24'b010100110010110000010000;
#10000;
	data_in <= 24'b010100100010101100001111;
#10000;
	data_in <= 24'b010100010010110000010010;
#10000;
	data_in <= 24'b010100100010110100010011;
#10000;
	data_in <= 24'b010100000010110000010100;
#10000;
	data_in <= 24'b010011110010101100010011;
#10000;
	data_in <= 24'b010011010010101100010100;
#10000;
	data_in <= 24'b010011100010110000010101;
#10000;
	data_in <= 24'b010101010010111000010010;
#10000;
	data_in <= 24'b010100110010111000010010;
#10000;
	data_in <= 24'b010100110010111000010100;
#10000;
	data_in <= 24'b010100110011000000010110;
#10000;
	data_in <= 24'b010100100010111000010110;
#10000;
	data_in <= 24'b010011010010101100010011;
#10000;
	data_in <= 24'b010011000010101000010011;
#10000;
	data_in <= 24'b010011000010101000010011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001001100001010000001101;
#10000;
	data_in <= 24'b001010000001011000001111;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100000001110100010101;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001010000001011000001111;
#10000;
	data_in <= 24'b001010010001011100010000;
#10000;
	data_in <= 24'b001010110001100100010010;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100010001111000010110;
#10000;
	data_in <= 24'b001100100001111100010111;
#10000;
	data_in <= 24'b001010100001100000010001;
#10000;
	data_in <= 24'b001010110001100100010010;
#10000;
	data_in <= 24'b001011010001101000010011;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001100110010000000011000;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001010110001100100010010;
#10000;
	data_in <= 24'b001011000001101000010011;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001011000001100100010010;
#10000;
	data_in <= 24'b001011010001101000010011;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001010110001100000010001;
#10000;
	data_in <= 24'b001011010001101000010011;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001101010010001000011011;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001011000001100100010010;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001110000010001100011011;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001011010001101000010011;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001101000010000100011001;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001101110010001000011010;
#10000;
	data_in <= 24'b001110000010001100011011;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001110110010011100011100;
#10000;
	data_in <= 24'b001111000010100000011101;
#10000;
	data_in <= 24'b001111010010100100011110;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b001101110010001000011010;
#10000;
	data_in <= 24'b001110000010001100011011;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011100011100;
#10000;
	data_in <= 24'b001111000010100000011101;
#10000;
	data_in <= 24'b001111010010100100011110;
#10000;
	data_in <= 24'b001111110010100100011110;
#10000;
	data_in <= 24'b001101110010001000011010;
#10000;
	data_in <= 24'b001110000010001100011011;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111000010100000011101;
#10000;
	data_in <= 24'b001111000010100000011101;
#10000;
	data_in <= 24'b001111110010100100011110;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b001110000010001100011011;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111010010100100011110;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111010010100100011110;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111000010100000011101;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111010010100100011110;
#10000;
	data_in <= 24'b001111100010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000000010101000011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010000110010110100100001;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010000010010100100011101;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010001100010111100100000;
#10000;
	data_in <= 24'b010010000011000100100010;
#10000;
	data_in <= 24'b010010010011000000100000;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010000100010101000011110;
#10000;
	data_in <= 24'b010000010010100100011101;
#10000;
	data_in <= 24'b010000100010101000011110;
#10000;
	data_in <= 24'b010001010010111000011111;
#10000;
	data_in <= 24'b010001110011000000100001;
#10000;
	data_in <= 24'b010010010011000000100000;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010010000010111000100000;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010001010010110100100001;
#10000;
	data_in <= 24'b010001010010110100100001;
#10000;
	data_in <= 24'b010001100010111000100010;
#10000;
	data_in <= 24'b010001100010111000100010;
#10000;
	data_in <= 24'b010010000010111000100000;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010001100010110000011110;
#10000;
	data_in <= 24'b010001100010110000011110;
#10000;
	data_in <= 24'b010001100010110000011110;
#10000;
	data_in <= 24'b010001110010110100011111;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010010010011000000100000;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010001100010110000011110;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010001100010110000011110;
#10000;
	data_in <= 24'b010001110010111000011110;
#10000;
	data_in <= 24'b010010010011000000100000;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010001000010101000011110;
#10000;
	data_in <= 24'b010001000010101000011100;
#10000;
	data_in <= 24'b010001000010101000011100;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010010000010111100011111;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010011100011010100100101;
#10000;
	data_in <= 24'b010011110011011000100110;
#10000;
	data_in <= 24'b010100000011011000100110;
#10000;
	data_in <= 24'b010100000011011000100110;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010010010011000000100000;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010011010011010000100100;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010010100011000100100001;
#10000;
	data_in <= 24'b010011000011001100100011;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011110011010100100101;
#10000;
	data_in <= 24'b010011110011010100100101;
#10000;
	data_in <= 24'b010011110011010100100101;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010010100011000000100000;
#10000;
	data_in <= 24'b010010110011000100100001;
#10000;
	data_in <= 24'b010011000011001000100010;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010100100011010100100111;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
	data_in <= 24'b010010100011000000100000;
#10000;
	data_in <= 24'b010010110011000100100001;
#10000;
	data_in <= 24'b010011000011001000100010;
#10000;
	data_in <= 24'b010011000011001000100010;
#10000;
	data_in <= 24'b010011000011001000100010;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010100010011010000100110;
#10000;
	data_in <= 24'b010100110011011000101000;
#10000;
	data_in <= 24'b010011000011001000100010;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011100011000100100010;
#10000;
	data_in <= 24'b010011110011001000100011;
#10000;
	data_in <= 24'b010100010011010000100110;
#10000;
	data_in <= 24'b010100110011011000101000;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010011010011001100100011;
#10000;
	data_in <= 24'b010011000011001000100010;
#10000;
	data_in <= 24'b010011010011000000100001;
#10000;
	data_in <= 24'b010011010011000000100001;
#10000;
	data_in <= 24'b010011110011001000100100;
#10000;
	data_in <= 24'b010100010011010000100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100010011011100100111;
#10000;
	data_in <= 24'b010100000011011000100110;
#10000;
	data_in <= 24'b010100000011011000100110;
#10000;
	data_in <= 24'b010100010011011100100111;
#10000;
	data_in <= 24'b010100100011011000100101;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010011100011001000100001;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010100110011100100101001;
#10000;
	data_in <= 24'b010100100011100000101000;
#10000;
	data_in <= 24'b010100010011011100100111;
#10000;
	data_in <= 24'b010100010011011100100111;
#10000;
	data_in <= 24'b010100100011011000100101;
#10000;
	data_in <= 24'b010011110011001100100010;
#10000;
	data_in <= 24'b010011010011000100100000;
#10000;
	data_in <= 24'b010011010011000100100000;
#10000;
	data_in <= 24'b010100010011011100100111;
#10000;
	data_in <= 24'b010100000011011000100110;
#10000;
	data_in <= 24'b010100010011010000100101;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100100011010000100011;
#10000;
	data_in <= 24'b010100100011010000100011;
#10000;
	data_in <= 24'b010100000011011000100110;
#10000;
	data_in <= 24'b010011100011010000100100;
#10000;
	data_in <= 24'b010100000011001100100100;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010101000011011100101000;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010101010011011100100110;
#10000;
	data_in <= 24'b010101000011011000100101;
#10000;
	data_in <= 24'b010101100011100100101010;
#10000;
	data_in <= 24'b010101000011011100101000;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100010011010000100101;
#10000;
	data_in <= 24'b010100100011001100100100;
#10000;
	data_in <= 24'b010100010011001100100010;
#10000;
	data_in <= 24'b010101100011100100101010;
#10000;
	data_in <= 24'b010101010011100000101001;
#10000;
	data_in <= 24'b010101000011011100101000;
#10000;
	data_in <= 24'b010101000011011100101000;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100000011001100100100;
#10000;
	data_in <= 24'b010100010011001000100011;
#10000;
	data_in <= 24'b010100100011001100100100;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100010011010000100101;
#10000;
	data_in <= 24'b010101000011010100100110;
#10000;
	data_in <= 24'b010101100011011100101000;
#10000;
	data_in <= 24'b010100010011010000100101;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100110011011000100111;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100000011001100100100;
#10000;
	data_in <= 24'b010101000011010100100110;
#10000;
	data_in <= 24'b010101110011100000101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100100011010000100001;
#10000;
	data_in <= 24'b010100100011010000100001;
#10000;
	data_in <= 24'b010101000011010100100000;
#10000;
	data_in <= 24'b010100110011010000011111;
#10000;
	data_in <= 24'b010100010011001000011101;
#10000;
	data_in <= 24'b010011110011000000011011;
#10000;
	data_in <= 24'b010100010011001000011011;
#10000;
	data_in <= 24'b010101000011010100011110;
#10000;
	data_in <= 24'b010011110011000100011110;
#10000;
	data_in <= 24'b010011110011000100011110;
#10000;
	data_in <= 24'b010100010011001000011101;
#10000;
	data_in <= 24'b010100010011001000011101;
#10000;
	data_in <= 24'b010100000011000100011100;
#10000;
	data_in <= 24'b010100000011000100011100;
#10000;
	data_in <= 24'b010100010011001000011101;
#10000;
	data_in <= 24'b010101000011010100011110;
#10000;
	data_in <= 24'b010100010011001100100000;
#10000;
	data_in <= 24'b010100000011001000011111;
#10000;
	data_in <= 24'b010100010011000100011110;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100110011001100100000;
#10000;
	data_in <= 24'b010100110011010000011111;
#10000;
	data_in <= 24'b010101000011010100100000;
#10000;
	data_in <= 24'b010101100011011100100010;
#10000;
	data_in <= 24'b010101010011011100100110;
#10000;
	data_in <= 24'b010100110011010100100010;
#10000;
	data_in <= 24'b010101000011010000100001;
#10000;
	data_in <= 24'b010101010011010100100010;
#10000;
	data_in <= 24'b010101110011011100100100;
#10000;
	data_in <= 24'b010101110011011100100100;
#10000;
	data_in <= 24'b010101110011011100100100;
#10000;
	data_in <= 24'b010110000011100000100101;
#10000;
	data_in <= 24'b010101100011100000100111;
#10000;
	data_in <= 24'b010100110011010100100100;
#10000;
	data_in <= 24'b010101010011010000100100;
#10000;
	data_in <= 24'b010101100011010100100101;
#10000;
	data_in <= 24'b010110000011011100100111;
#10000;
	data_in <= 24'b010110010011100000101000;
#10000;
	data_in <= 24'b010110100011100000101000;
#10000;
	data_in <= 24'b010110100011100100101001;
#10000;
	data_in <= 24'b010101000011011000100101;
#10000;
	data_in <= 24'b010100110011010100100100;
#10000;
	data_in <= 24'b010101010011010000100100;
#10000;
	data_in <= 24'b010101110011011000100110;
#10000;
	data_in <= 24'b010110100011100100101001;
#10000;
	data_in <= 24'b010110110011101000101010;
#10000;
	data_in <= 24'b010111000011101000101010;
#10000;
	data_in <= 24'b010111000011101100101011;
#10000;
	data_in <= 24'b010101000011010100100110;
#10000;
	data_in <= 24'b010101000011010100100110;
#10000;
	data_in <= 24'b010101100011010100100110;
#10000;
	data_in <= 24'b010110010011100000101001;
#10000;
	data_in <= 24'b010110100011100100101010;
#10000;
	data_in <= 24'b010110110011101000101011;
#10000;
	data_in <= 24'b010111010011101000101100;
#10000;
	data_in <= 24'b010111100011110100101110;
#10000;
	data_in <= 24'b010101000011010100100110;
#10000;
	data_in <= 24'b010101000011010100100110;
#10000;
	data_in <= 24'b010101110011011000100111;
#10000;
	data_in <= 24'b010110000011011100101000;
#10000;
	data_in <= 24'b010110010011100000101001;
#10000;
	data_in <= 24'b010110010011100000101000;
#10000;
	data_in <= 24'b010110110011100000101010;
#10000;
	data_in <= 24'b010111000011101100101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100110011001000011110;
#10000;
	data_in <= 24'b010110100011100100100101;
#10000;
	data_in <= 24'b010111010011110000101000;
#10000;
	data_in <= 24'b010110100011100100100101;
#10000;
	data_in <= 24'b010101110011010100011110;
#10000;
	data_in <= 24'b010101010011001100011100;
#10000;
	data_in <= 24'b010101000011001000011011;
#10000;
	data_in <= 24'b010100110011000100011010;
#10000;
	data_in <= 24'b010100110011001000011110;
#10000;
	data_in <= 24'b010101010011010000100000;
#10000;
	data_in <= 24'b010101100011010100100001;
#10000;
	data_in <= 24'b010100110011001000011110;
#10000;
	data_in <= 24'b010101010011001100011100;
#10000;
	data_in <= 24'b010110010011011100100000;
#10000;
	data_in <= 24'b010110110011100100100010;
#10000;
	data_in <= 24'b010111000011101000100011;
#10000;
	data_in <= 24'b010100010011000100011110;
#10000;
	data_in <= 24'b010100100011001000011111;
#10000;
	data_in <= 24'b010100110011001000011110;
#10000;
	data_in <= 24'b010100110011001000011110;
#10000;
	data_in <= 24'b010101100011011000011111;
#10000;
	data_in <= 24'b010110100011101000100011;
#10000;
	data_in <= 24'b010111010011101100100011;
#10000;
	data_in <= 24'b010110100011100000100000;
#10000;
	data_in <= 24'b010101100011011000100011;
#10000;
	data_in <= 24'b010101100011011000100011;
#10000;
	data_in <= 24'b010101110011011000100011;
#10000;
	data_in <= 24'b010110000011011100100011;
#10000;
	data_in <= 24'b010110110011101000100110;
#10000;
	data_in <= 24'b010111110011111100101000;
#10000;
	data_in <= 24'b011000000011111000100110;
#10000;
	data_in <= 24'b010111010011101100100011;
#10000;
	data_in <= 24'b010111000011101100101011;
#10000;
	data_in <= 24'b010110100011110000101001;
#10000;
	data_in <= 24'b010110110011101100101000;
#10000;
	data_in <= 24'b010110110011110000100111;
#10000;
	data_in <= 24'b010111100011110100101001;
#10000;
	data_in <= 24'b011000100100001000101011;
#10000;
	data_in <= 24'b011010000100011000101110;
#10000;
	data_in <= 24'b011010100100100000110000;
#10000;
	data_in <= 24'b010110100011110000101011;
#10000;
	data_in <= 24'b010111000011111000101101;
#10000;
	data_in <= 24'b011000000011111100101111;
#10000;
	data_in <= 24'b011000000100000000101101;
#10000;
	data_in <= 24'b011000000011111100101011;
#10000;
	data_in <= 24'b011000100100001000101011;
#10000;
	data_in <= 24'b011001110100010100101110;
#10000;
	data_in <= 24'b011010100100100000110000;
#10000;
	data_in <= 24'b010110000011100100101010;
#10000;
	data_in <= 24'b010110100011111000101101;
#10000;
	data_in <= 24'b011000010100001100110010;
#10000;
	data_in <= 24'b011000010100001100110000;
#10000;
	data_in <= 24'b011000010100001000101101;
#10000;
	data_in <= 24'b010111100011111100101000;
#10000;
	data_in <= 24'b010111110011111100101000;
#10000;
	data_in <= 24'b011000000100000100101000;
#10000;
	data_in <= 24'b010110110011110000101101;
#10000;
	data_in <= 24'b010111100100000000101111;
#10000;
	data_in <= 24'b011000100100000100110001;
#10000;
	data_in <= 24'b011000010100000000110000;
#10000;
	data_in <= 24'b010111110011111000101011;
#10000;
	data_in <= 24'b010111100011110100101001;
#10000;
	data_in <= 24'b011000100100000000101001;
#10000;
	data_in <= 24'b011001010100001100101100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010101110011010100011110;
#10000;
	data_in <= 24'b010110110011100100100010;
#10000;
	data_in <= 24'b010111100011110100101001;
#10000;
	data_in <= 24'b011000000011111100101011;
#10000;
	data_in <= 24'b011000000011111100101100;
#10000;
	data_in <= 24'b011000000011111100101100;
#10000;
	data_in <= 24'b011000010100000100101110;
#10000;
	data_in <= 24'b011000100100001000101111;
#10000;
	data_in <= 24'b010110000011011000011111;
#10000;
	data_in <= 24'b010111000011101000100011;
#10000;
	data_in <= 24'b010111110011111000101010;
#10000;
	data_in <= 24'b011000000011111100101011;
#10000;
	data_in <= 24'b010111110011111000101011;
#10000;
	data_in <= 24'b010111100011110100101010;
#10000;
	data_in <= 24'b010111110011111100101100;
#10000;
	data_in <= 24'b011000110100001000101111;
#10000;
	data_in <= 24'b010111010011101100100011;
#10000;
	data_in <= 24'b011000010011111100100111;
#10000;
	data_in <= 24'b011001010100001100101100;
#10000;
	data_in <= 24'b011001000100001000101011;
#10000;
	data_in <= 24'b010111100011110100101001;
#10000;
	data_in <= 24'b010111000011101100100111;
#10000;
	data_in <= 24'b010111100011110100101001;
#10000;
	data_in <= 24'b011000010100000000101100;
#10000;
	data_in <= 24'b011001010100001100101011;
#10000;
	data_in <= 24'b011001110100010100101101;
#10000;
	data_in <= 24'b011010000100011000101111;
#10000;
	data_in <= 24'b011001010100001100101100;
#10000;
	data_in <= 24'b010111100011110100101001;
#10000;
	data_in <= 24'b010110100011100100100101;
#10000;
	data_in <= 24'b010110110011101000100110;
#10000;
	data_in <= 24'b010111010011110000101000;
#10000;
	data_in <= 24'b011010000100011000101110;
#10000;
	data_in <= 24'b011010000100011000101110;
#10000;
	data_in <= 24'b011001100100010000101100;
#10000;
	data_in <= 24'b011000100100000000101000;
#10000;
	data_in <= 24'b010111100011110000100101;
#10000;
	data_in <= 24'b010110110011100100100010;
#10000;
	data_in <= 24'b010110100011100000100001;
#10000;
	data_in <= 24'b010110110011100000100100;
#10000;
	data_in <= 24'b011001100100010000101100;
#10000;
	data_in <= 24'b011001010100001100101011;
#10000;
	data_in <= 24'b011000100100000000101000;
#10000;
	data_in <= 24'b010111110011110100100101;
#10000;
	data_in <= 24'b010110110011100100100010;
#10000;
	data_in <= 24'b010110100011100000100001;
#10000;
	data_in <= 24'b010110010011011100100000;
#10000;
	data_in <= 24'b010110100011100000100001;
#10000;
	data_in <= 24'b011001100100010100101011;
#10000;
	data_in <= 24'b011001010100010000101010;
#10000;
	data_in <= 24'b011001010100001000101000;
#10000;
	data_in <= 24'b011000010011111000100100;
#10000;
	data_in <= 24'b010111010011100100100001;
#10000;
	data_in <= 24'b010111000011100000100000;
#10000;
	data_in <= 24'b010111010011100000100010;
#10000;
	data_in <= 24'b010111110011101000100100;
#10000;
	data_in <= 24'b011010000100011000101110;
#10000;
	data_in <= 24'b011010000100011000101110;
#10000;
	data_in <= 24'b011010000100010000101100;
#10000;
	data_in <= 24'b011000110011111100100111;
#10000;
	data_in <= 24'b010111100011101000100010;
#10000;
	data_in <= 24'b010110100011100000100000;
#10000;
	data_in <= 24'b010111010011101100100100;
#10000;
	data_in <= 24'b011000000011111000100111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011001010100010000110001;
#10000;
	data_in <= 24'b011000010011110100101011;
#10000;
	data_in <= 24'b010111000011100000100110;
#10000;
	data_in <= 24'b010111100011101000101000;
#10000;
	data_in <= 24'b011000100011111000101100;
#10000;
	data_in <= 24'b011000100011111000101100;
#10000;
	data_in <= 24'b010111100011100100100101;
#10000;
	data_in <= 24'b010110010011010000100000;
#10000;
	data_in <= 24'b011001010100000100101111;
#10000;
	data_in <= 24'b011000010011110100101011;
#10000;
	data_in <= 24'b010111100011101000101000;
#10000;
	data_in <= 24'b010111110011101100101001;
#10000;
	data_in <= 24'b011000000011110000101010;
#10000;
	data_in <= 24'b010111110011110000101000;
#10000;
	data_in <= 24'b010111100011100100100101;
#10000;
	data_in <= 24'b010111000011011100100001;
#10000;
	data_in <= 24'b011000100011111000101100;
#10000;
	data_in <= 24'b011000100011111000101100;
#10000;
	data_in <= 24'b011000010011110100101011;
#10000;
	data_in <= 24'b011000010011110100101011;
#10000;
	data_in <= 24'b011000010011110000101000;
#10000;
	data_in <= 24'b010111100011100100100101;
#10000;
	data_in <= 24'b010111010011100000100100;
#10000;
	data_in <= 24'b010111100011100100100011;
#10000;
	data_in <= 24'b011000000011110000101010;
#10000;
	data_in <= 24'b011000010011110100101011;
#10000;
	data_in <= 24'b011000100011111000101100;
#10000;
	data_in <= 24'b011000100011111000101100;
#10000;
	data_in <= 24'b011000010011110000101000;
#10000;
	data_in <= 24'b010111010011100000100100;
#10000;
	data_in <= 24'b010111000011011100100001;
#10000;
	data_in <= 24'b010111010011100000100010;
#10000;
	data_in <= 24'b010111000011100000100110;
#10000;
	data_in <= 24'b010111010011100100100111;
#10000;
	data_in <= 24'b010111110011101100101001;
#10000;
	data_in <= 24'b011000010011110100101011;
#10000;
	data_in <= 24'b010111110011110000101000;
#10000;
	data_in <= 24'b010111000011100100100101;
#10000;
	data_in <= 24'b010111010011100000100010;
#10000;
	data_in <= 24'b010111010011100000100010;
#10000;
	data_in <= 24'b010110100011011000100100;
#10000;
	data_in <= 24'b010110100011011000100100;
#10000;
	data_in <= 24'b010111000011100000100110;
#10000;
	data_in <= 24'b010111100011101000101000;
#10000;
	data_in <= 24'b010111110011110000101000;
#10000;
	data_in <= 24'b010111100011101100100111;
#10000;
	data_in <= 24'b010111100011100100100011;
#10000;
	data_in <= 24'b010111100011100100100011;
#10000;
	data_in <= 24'b010111110011101100101001;
#10000;
	data_in <= 24'b010111010011100100100111;
#10000;
	data_in <= 24'b010111010011100100100111;
#10000;
	data_in <= 24'b010111100011101000101000;
#10000;
	data_in <= 24'b010111110011110000101000;
#10000;
	data_in <= 24'b010111100011101100100111;
#10000;
	data_in <= 24'b010111100011110000100101;
#10000;
	data_in <= 24'b010111110011110100100110;
#10000;
	data_in <= 24'b011001010100001000101110;
#10000;
	data_in <= 24'b011000110100000000101100;
#10000;
	data_in <= 24'b011000010011111000101010;
#10000;
	data_in <= 24'b011000000011110100101001;
#10000;
	data_in <= 24'b010111100011101100100111;
#10000;
	data_in <= 24'b010111100011110000100101;
#10000;
	data_in <= 24'b010111100011110000100101;
#10000;
	data_in <= 24'b011000000011111000100111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010110110011010000011110;
#10000;
	data_in <= 24'b010101010010111100010111;
#10000;
	data_in <= 24'b010111010011010100011100;
#10000;
	data_in <= 24'b010110010011000100010101;
#10000;
	data_in <= 24'b011110100100111100110100;
#10000;
	data_in <= 24'b100001000101101000111101;
#10000;
	data_in <= 24'b010110010010110100010000;
#10000;
	data_in <= 24'b010110110011001000010010;
#10000;
	data_in <= 24'b011000010011101100100011;
#10000;
	data_in <= 24'b010111100011100100011111;
#10000;
	data_in <= 24'b011001000011101100100010;
#10000;
	data_in <= 24'b011000010011100100011101;
#10000;
	data_in <= 24'b011011110100010100101000;
#10000;
	data_in <= 24'b011100110100100100101100;
#10000;
	data_in <= 24'b011000110011011100011000;
#10000;
	data_in <= 24'b011000010011100000011000;
#10000;
	data_in <= 24'b010111110011100100100001;
#10000;
	data_in <= 24'b010111010011100000011110;
#10000;
	data_in <= 24'b010111110011011000011101;
#10000;
	data_in <= 24'b011000010011100100011101;
#10000;
	data_in <= 24'b010111110011010100011000;
#10000;
	data_in <= 24'b011000000011011100010111;
#10000;
	data_in <= 24'b011001100011101000011011;
#10000;
	data_in <= 24'b010111100011010100010101;
#10000;
	data_in <= 24'b010111110011100100100001;
#10000;
	data_in <= 24'b010111010011100000011110;
#10000;
	data_in <= 24'b010110110011001100011010;
#10000;
	data_in <= 24'b011000000011100000011100;
#10000;
	data_in <= 24'b011000000011011000011001;
#10000;
	data_in <= 24'b010111110011011000010110;
#10000;
	data_in <= 24'b011010000011110000011101;
#10000;
	data_in <= 24'b010111010011010000010100;
#10000;
	data_in <= 24'b011000000011101000100010;
#10000;
	data_in <= 24'b010111010011100000011110;
#10000;
	data_in <= 24'b010111000011010000011011;
#10000;
	data_in <= 24'b010111010011011000011010;
#10000;
	data_in <= 24'b011000100011101000011101;
#10000;
	data_in <= 24'b011000100011101000011101;
#10000;
	data_in <= 24'b011000010011100000011000;
#10000;
	data_in <= 24'b010111110011011000010110;
#10000;
	data_in <= 24'b011000000011101000100010;
#10000;
	data_in <= 24'b010111010011011100011111;
#10000;
	data_in <= 24'b010111100011011000011101;
#10000;
	data_in <= 24'b010110100011001100010111;
#10000;
	data_in <= 24'b010111110011011100011010;
#10000;
	data_in <= 24'b011000000011100000011011;
#10000;
	data_in <= 24'b010110100011000100010001;
#10000;
	data_in <= 24'b011000000011011100010111;
#10000;
	data_in <= 24'b011000110011111100100111;
#10000;
	data_in <= 24'b011000000011110000100100;
#10000;
	data_in <= 24'b011000000011101100100001;
#10000;
	data_in <= 24'b010111100011100100011101;
#10000;
	data_in <= 24'b011000000011101000011100;
#10000;
	data_in <= 24'b010111110011100100011011;
#10000;
	data_in <= 24'b010111010011011000010110;
#10000;
	data_in <= 24'b011000000011100100011001;
#10000;
	data_in <= 24'b011001100100001000101010;
#10000;
	data_in <= 24'b011000000011110000100100;
#10000;
	data_in <= 24'b010111100011100100011111;
#10000;
	data_in <= 24'b011000100011110100100011;
#10000;
	data_in <= 24'b011000010011101000011110;
#10000;
	data_in <= 24'b010111110011100000011100;
#10000;
	data_in <= 24'b011000010011101100011101;
#10000;
	data_in <= 24'b010111000011010000010111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010111010011001100010110;
#10000;
	data_in <= 24'b010110110011001100010110;
#10000;
	data_in <= 24'b010110100011001000010101;
#10000;
	data_in <= 24'b010110010011000100010100;
#10000;
	data_in <= 24'b010101110010111100010010;
#10000;
	data_in <= 24'b010101110010111100010010;
#10000;
	data_in <= 24'b010110010011000100010100;
#10000;
	data_in <= 24'b010110100011010000010110;
#10000;
	data_in <= 24'b010111000011010000010111;
#10000;
	data_in <= 24'b010110110011001100010110;
#10000;
	data_in <= 24'b010110010011000100010100;
#10000;
	data_in <= 24'b010110000011000000010011;
#10000;
	data_in <= 24'b010110000011000000010011;
#10000;
	data_in <= 24'b010110000011000000010011;
#10000;
	data_in <= 24'b010101110011000100010011;
#10000;
	data_in <= 24'b010101110011000100010011;
#10000;
	data_in <= 24'b010111010011011000010110;
#10000;
	data_in <= 24'b010110100011010000010100;
#10000;
	data_in <= 24'b010110000011001000010010;
#10000;
	data_in <= 24'b010110000011001000010010;
#10000;
	data_in <= 24'b010110000011001000010010;
#10000;
	data_in <= 24'b010110000011001000010010;
#10000;
	data_in <= 24'b010101110011000100010001;
#10000;
	data_in <= 24'b010101010010111100001111;
#10000;
	data_in <= 24'b010110110011010000010100;
#10000;
	data_in <= 24'b010110010011001100010011;
#10000;
	data_in <= 24'b010110000011001000010010;
#10000;
	data_in <= 24'b010110000011001000010010;
#10000;
	data_in <= 24'b010110000011001000010010;
#10000;
	data_in <= 24'b010110000011001000010010;
#10000;
	data_in <= 24'b010101110011000100010001;
#10000;
	data_in <= 24'b010101100011000000010000;
#10000;
	data_in <= 24'b010110010011001000010010;
#10000;
	data_in <= 24'b010110100011001100010011;
#10000;
	data_in <= 24'b010110110011010000010100;
#10000;
	data_in <= 24'b010110100011001100010011;
#10000;
	data_in <= 24'b010110010011001000010010;
#10000;
	data_in <= 24'b010110010011001000010010;
#10000;
	data_in <= 24'b010110010011001000010010;
#10000;
	data_in <= 24'b010110010011001000010010;
#10000;
	data_in <= 24'b010110010011001000010010;
#10000;
	data_in <= 24'b010110110011010000010100;
#10000;
	data_in <= 24'b010111000011010100010101;
#10000;
	data_in <= 24'b010110110011010000010100;
#10000;
	data_in <= 24'b010110100011001100010011;
#10000;
	data_in <= 24'b010110010011001000010010;
#10000;
	data_in <= 24'b010110100011001100010011;
#10000;
	data_in <= 24'b010110110011010000010100;
#10000;
	data_in <= 24'b010111010011011000010110;
#10000;
	data_in <= 24'b010111010011011000010110;
#10000;
	data_in <= 24'b010111110011011000010110;
#10000;
	data_in <= 24'b010111100011010100010101;
#10000;
	data_in <= 24'b010111100011010100010101;
#10000;
	data_in <= 24'b010111010011010000010100;
#10000;
	data_in <= 24'b010111100011010100010101;
#10000;
	data_in <= 24'b010111100011010100010101;
#10000;
	data_in <= 24'b011000000011100100011001;
#10000;
	data_in <= 24'b010111100011011100010111;
#10000;
	data_in <= 24'b010111110011011000010110;
#10000;
	data_in <= 24'b010111100011010100010101;
#10000;
	data_in <= 24'b010111110011011000010110;
#10000;
	data_in <= 24'b010111110011011000010110;
#10000;
	data_in <= 24'b010111110011011000010110;
#10000;
	data_in <= 24'b010111000011010100010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010101010010111100010001;
#10000;
	data_in <= 24'b010101000011000000010010;
#10000;
	data_in <= 24'b010101000010111100010011;
#10000;
	data_in <= 24'b010100000010110100010011;
#10000;
	data_in <= 24'b010011100010101000010010;
#10000;
	data_in <= 24'b010011000010101000010010;
#10000;
	data_in <= 24'b010011100010110000010100;
#10000;
	data_in <= 24'b010011110011000000010111;
#10000;
	data_in <= 24'b010101000011000000010010;
#10000;
	data_in <= 24'b010101000011000000010010;
#10000;
	data_in <= 24'b010100100011000000010011;
#10000;
	data_in <= 24'b010100100011000000010011;
#10000;
	data_in <= 24'b010100000010111100010101;
#10000;
	data_in <= 24'b010100010010111100010111;
#10000;
	data_in <= 24'b010100010011001000011001;
#10000;
	data_in <= 24'b010100100011001100011010;
#10000;
	data_in <= 24'b010101010011000100010011;
#10000;
	data_in <= 24'b010101010011000100010011;
#10000;
	data_in <= 24'b010100110011000100010100;
#10000;
	data_in <= 24'b010101010011001100010110;
#10000;
	data_in <= 24'b010101010011010000011010;
#10000;
	data_in <= 24'b010101110011011000011100;
#10000;
	data_in <= 24'b010101010011011000011101;
#10000;
	data_in <= 24'b010101010011011000011101;
#10000;
	data_in <= 24'b010110010011001100010101;
#10000;
	data_in <= 24'b010101110011001100010101;
#10000;
	data_in <= 24'b010110000011001100010111;
#10000;
	data_in <= 24'b010110000011011000011001;
#10000;
	data_in <= 24'b010110010011011000011100;
#10000;
	data_in <= 24'b010110000011011100011101;
#10000;
	data_in <= 24'b010101110011010100011101;
#10000;
	data_in <= 24'b010101010011011000011101;
#10000;
	data_in <= 24'b010110110011001100010110;
#10000;
	data_in <= 24'b010111000011011000011000;
#10000;
	data_in <= 24'b010111010011011000011010;
#10000;
	data_in <= 24'b010110110011011000011010;
#10000;
	data_in <= 24'b010110110011011000011100;
#10000;
	data_in <= 24'b010101110011010000011010;
#10000;
	data_in <= 24'b010101100011001000011010;
#10000;
	data_in <= 24'b010101000011001000011010;
#10000;
	data_in <= 24'b010111000011010000010111;
#10000;
	data_in <= 24'b010111010011010100011000;
#10000;
	data_in <= 24'b010111110011011100011011;
#10000;
	data_in <= 24'b010111010011011000011010;
#10000;
	data_in <= 24'b010111000011010000011011;
#10000;
	data_in <= 24'b010101110011001000011000;
#10000;
	data_in <= 24'b010101100011000000011000;
#10000;
	data_in <= 24'b010100110010111100010111;
#10000;
	data_in <= 24'b010111100011010000010111;
#10000;
	data_in <= 24'b010111000011010000010111;
#10000;
	data_in <= 24'b010111010011010100011001;
#10000;
	data_in <= 24'b010111010011010100011001;
#10000;
	data_in <= 24'b010111010011010000011011;
#10000;
	data_in <= 24'b010110110011001000011011;
#10000;
	data_in <= 24'b010110010011000000011001;
#10000;
	data_in <= 24'b010101010010111100010111;
#10000;
	data_in <= 24'b010111100011010000010111;
#10000;
	data_in <= 24'b010110110011001100010110;
#10000;
	data_in <= 24'b010110110011001100010111;
#10000;
	data_in <= 24'b010111000011010000011000;
#10000;
	data_in <= 24'b010111100011010100011100;
#10000;
	data_in <= 24'b010111100011010100011100;
#10000;
	data_in <= 24'b010110110011001000011011;
#10000;
	data_in <= 24'b010110000011000000010111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001011000001100100010010;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001101100010001100011011;
#10000;
	data_in <= 24'b001101110010010000011100;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001011010001101000010011;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001101010010001000011010;
#10000;
	data_in <= 24'b001101110010010000011100;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001101010010001000011011;
#10000;
	data_in <= 24'b001101110010010000011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001101010010001000011011;
#10000;
	data_in <= 24'b001101110010010000011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001101100010001100011100;
#10000;
	data_in <= 24'b001110000010010100011110;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001011100001101100010100;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001101100010001100011100;
#10000;
	data_in <= 24'b001110000010010100011110;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001011110001110000010101;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001101010010001000011011;
#10000;
	data_in <= 24'b001101110010010000011101;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100000001110100010110;
#10000;
	data_in <= 24'b001100010001111000010111;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001101000010000100011010;
#10000;
	data_in <= 24'b001101100010001100011100;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010000110010110100100001;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010000110010110100100001;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111110010101100100000;
#10000;
	data_in <= 24'b010000010010110100100010;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000010010110100100010;
#10000;
	data_in <= 24'b010000110010111100100100;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001100011000000100101;
#10000;
	data_in <= 24'b010001100011000000100101;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001010010111100100011;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001110010111100100011;
#10000;
	data_in <= 24'b001111110010100000100000;
#10000;
	data_in <= 24'b010000000010100100100001;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001100010110100100011;
#10000;
	data_in <= 24'b010001100010111000100010;
#10000;
	data_in <= 24'b001111100010011100011111;
#10000;
	data_in <= 24'b001111100010011100011111;
#10000;
	data_in <= 24'b001111110010100100011110;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000010010101100100000;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010001010010110000100010;
#10000;
	data_in <= 24'b010001100010111000100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010001100010110000100000;
#10000;
	data_in <= 24'b010001010010101100011101;
#10000;
	data_in <= 24'b010001100010110000011110;
#10000;
	data_in <= 24'b010001110010110100011111;
#10000;
	data_in <= 24'b010010000010111000100000;
#10000;
	data_in <= 24'b010010000010111000100000;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010011010011001100100101;
#10000;
	data_in <= 24'b010010010010111100100011;
#10000;
	data_in <= 24'b010010000010111000100000;
#10000;
	data_in <= 24'b010010000010111000100000;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010011010011001100100101;
#10000;
	data_in <= 24'b010010110011000100100101;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010010110011000100100101;
#10000;
	data_in <= 24'b010010110011000100100011;
#10000;
	data_in <= 24'b010010110011000100100011;
#10000;
	data_in <= 24'b010010110011000100100011;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010010110011000100100011;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010010010010111100100011;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010010100011000000100010;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010010000010111000100010;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010010010111100100001;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010010000010111000100010;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010010010010111000100000;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010101000011100100101011;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010101010011101000101100;
#10000;
	data_in <= 24'b010101010011101000101100;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010101010011101000101100;
#10000;
	data_in <= 24'b010101100011101100101101;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010101000011100100101011;
#10000;
	data_in <= 24'b010101100011101100101101;
#10000;
	data_in <= 24'b010110000011110100101111;
#10000;
	data_in <= 24'b010110010011111000110000;
#10000;
	data_in <= 24'b010110100011111100110001;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010101010011101000101100;
#10000;
	data_in <= 24'b010110010011111000110000;
#10000;
	data_in <= 24'b010110100011111100110001;
#10000;
	data_in <= 24'b010110100011111100110001;
#10000;
	data_in <= 24'b010110010011111000110000;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010101000011100100101011;
#10000;
	data_in <= 24'b010101100011101100101101;
#10000;
	data_in <= 24'b010101110011110000101110;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010110100011110100101111;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010100110011100000101010;
#10000;
	data_in <= 24'b010110000011101100101101;
#10000;
	data_in <= 24'b010111000011111100110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100000011001100100100;
#10000;
	data_in <= 24'b010011110011001000100011;
#10000;
	data_in <= 24'b010011110011001000100011;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010101010011011000100111;
#10000;
	data_in <= 24'b010101000011010100100110;
#10000;
	data_in <= 24'b010100110011010100100100;
#10000;
	data_in <= 24'b010100110011010100100100;
#10000;
	data_in <= 24'b010101000011011100101000;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100000011001100100100;
#10000;
	data_in <= 24'b010100010011010000100101;
#10000;
	data_in <= 24'b010100110011010000100101;
#10000;
	data_in <= 24'b010100100011001100100100;
#10000;
	data_in <= 24'b010100100011010000100011;
#10000;
	data_in <= 24'b010100100011010000100011;
#10000;
	data_in <= 24'b010101010011100000101001;
#10000;
	data_in <= 24'b010100100011010100100110;
#10000;
	data_in <= 24'b010100010011010000100101;
#10000;
	data_in <= 24'b010100010011010000100101;
#10000;
	data_in <= 24'b010100110011010000100101;
#10000;
	data_in <= 24'b010101000011010100100110;
#10000;
	data_in <= 24'b010101010011011100100110;
#10000;
	data_in <= 24'b010101100011100000100111;
#10000;
	data_in <= 24'b010101110011101000101011;
#10000;
	data_in <= 24'b010101010011100000101001;
#10000;
	data_in <= 24'b010101000011011100101000;
#10000;
	data_in <= 24'b010101000011011100101000;
#10000;
	data_in <= 24'b010101110011100000101001;
#10000;
	data_in <= 24'b010101110011100000101001;
#10000;
	data_in <= 24'b010110010011101100101010;
#10000;
	data_in <= 24'b010110100011110000101011;
#10000;
	data_in <= 24'b010110110011111000101111;
#10000;
	data_in <= 24'b010110100011110100101110;
#10000;
	data_in <= 24'b010110010011110000101101;
#10000;
	data_in <= 24'b010110100011110100101110;
#10000;
	data_in <= 24'b010110110011110000101101;
#10000;
	data_in <= 24'b010110100011101100101100;
#10000;
	data_in <= 24'b010110100011110000101011;
#10000;
	data_in <= 24'b010110110011110100101100;
#10000;
	data_in <= 24'b010110110011111000101111;
#10000;
	data_in <= 24'b010110110011111000101111;
#10000;
	data_in <= 24'b010110110011111000101111;
#10000;
	data_in <= 24'b010111010100000000110001;
#10000;
	data_in <= 24'b010111100011111100110000;
#10000;
	data_in <= 24'b010111010011111000101111;
#10000;
	data_in <= 24'b010111010011111100101110;
#10000;
	data_in <= 24'b010111100100000000101111;
#10000;
	data_in <= 24'b010110000011101100101100;
#10000;
	data_in <= 24'b010110000011101100101100;
#10000;
	data_in <= 24'b010110100011110100101110;
#10000;
	data_in <= 24'b010111000011111100110000;
#10000;
	data_in <= 24'b010111100011111100110000;
#10000;
	data_in <= 24'b010111010011111000101111;
#10000;
	data_in <= 24'b010111100100000000101111;
#10000;
	data_in <= 24'b011000000100001000110001;
#10000;
	data_in <= 24'b010110010011110000101101;
#10000;
	data_in <= 24'b010110010011110000101101;
#10000;
	data_in <= 24'b010110100011110100101110;
#10000;
	data_in <= 24'b010110110011111000101111;
#10000;
	data_in <= 24'b010111000011110100101110;
#10000;
	data_in <= 24'b010110110011110000101101;
#10000;
	data_in <= 24'b010111000011111000101101;
#10000;
	data_in <= 24'b010111010011111100101110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010101110011011000100110;
#10000;
	data_in <= 24'b010101100011010100100101;
#10000;
	data_in <= 24'b010101110011010100100101;
#10000;
	data_in <= 24'b010110010011011100100111;
#10000;
	data_in <= 24'b010110100011100000101000;
#10000;
	data_in <= 24'b010111000011101100101000;
#10000;
	data_in <= 24'b010111100011110000101100;
#10000;
	data_in <= 24'b011000010100000000101101;
#10000;
	data_in <= 24'b010101110011011000100110;
#10000;
	data_in <= 24'b010101010011010000100100;
#10000;
	data_in <= 24'b010101100011010000100100;
#10000;
	data_in <= 24'b010110000011011000100110;
#10000;
	data_in <= 24'b010110100011100100100110;
#10000;
	data_in <= 24'b010110110011101000100111;
#10000;
	data_in <= 24'b010111100011110100101010;
#10000;
	data_in <= 24'b011000000011111100101100;
#10000;
	data_in <= 24'b010110010011100000101000;
#10000;
	data_in <= 24'b010110000011011100100111;
#10000;
	data_in <= 24'b010110010011011100100111;
#10000;
	data_in <= 24'b010110100011100000101000;
#10000;
	data_in <= 24'b010110110011101000100111;
#10000;
	data_in <= 24'b010111010011110000101001;
#10000;
	data_in <= 24'b010111110011111000101011;
#10000;
	data_in <= 24'b011000100100000100101110;
#10000;
	data_in <= 24'b010111010011110000101100;
#10000;
	data_in <= 24'b010111000011101100101011;
#10000;
	data_in <= 24'b010111000011101000101010;
#10000;
	data_in <= 24'b010111010011101100101011;
#10000;
	data_in <= 24'b010111010011110000101001;
#10000;
	data_in <= 24'b010111100011110100101010;
#10000;
	data_in <= 24'b010111110011111000101011;
#10000;
	data_in <= 24'b011000010100000000101101;
#10000;
	data_in <= 24'b010111110011111000101110;
#10000;
	data_in <= 24'b010111100011110100101101;
#10000;
	data_in <= 24'b010111100011110000101100;
#10000;
	data_in <= 24'b010111100011110000101100;
#10000;
	data_in <= 24'b010111100011110100101010;
#10000;
	data_in <= 24'b010111010011110000101001;
#10000;
	data_in <= 24'b010111010011110000101001;
#10000;
	data_in <= 24'b010111110011111000101010;
#10000;
	data_in <= 24'b011000100100000100110001;
#10000;
	data_in <= 24'b011000010100000000110000;
#10000;
	data_in <= 24'b011000100100000000110000;
#10000;
	data_in <= 24'b011000110100000100110001;
#10000;
	data_in <= 24'b011000110100001000101111;
#10000;
	data_in <= 24'b011000010100000000101101;
#10000;
	data_in <= 24'b011000000011111100101100;
#10000;
	data_in <= 24'b011000010100000000101100;
#10000;
	data_in <= 24'b011001010100010000110100;
#10000;
	data_in <= 24'b011001010100010000110100;
#10000;
	data_in <= 24'b011001110100010100110101;
#10000;
	data_in <= 24'b011010100100100000111000;
#10000;
	data_in <= 24'b011010100100100100110110;
#10000;
	data_in <= 24'b011010010100100000110101;
#10000;
	data_in <= 24'b011010000100011100110100;
#10000;
	data_in <= 24'b011010000100011100110011;
#10000;
	data_in <= 24'b011001100100010100110101;
#10000;
	data_in <= 24'b011001100100010100110101;
#10000;
	data_in <= 24'b011010100100100000111000;
#10000;
	data_in <= 24'b011011100100110000111100;
#10000;
	data_in <= 24'b011011110100111000111011;
#10000;
	data_in <= 24'b011011100100110100111010;
#10000;
	data_in <= 24'b011011100100110100111010;
#10000;
	data_in <= 24'b011011100100110100111001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011000110100001000110010;
#10000;
	data_in <= 24'b010111110011111000101110;
#10000;
	data_in <= 24'b011001000100001000110010;
#10000;
	data_in <= 24'b011000110100000100110001;
#10000;
	data_in <= 24'b011010100100011000110110;
#10000;
	data_in <= 24'b011001010100000100101111;
#10000;
	data_in <= 24'b011010100100010000110010;
#10000;
	data_in <= 24'b011010100100010000110010;
#10000;
	data_in <= 24'b011000110100001000101111;
#10000;
	data_in <= 24'b011000010100000000101101;
#10000;
	data_in <= 24'b011010100100011000110100;
#10000;
	data_in <= 24'b011000110011111100101101;
#10000;
	data_in <= 24'b011010010100001100110001;
#10000;
	data_in <= 24'b011001100100000000101110;
#10000;
	data_in <= 24'b011100110100101100111001;
#10000;
	data_in <= 24'b011100100100101000111000;
#10000;
	data_in <= 24'b011000110100001000101110;
#10000;
	data_in <= 24'b010111110011111000101010;
#10000;
	data_in <= 24'b011010010100011000110010;
#10000;
	data_in <= 24'b011001100100001100101111;
#10000;
	data_in <= 24'b011011000100011100110011;
#10000;
	data_in <= 24'b011011010100100000110100;
#10000;
	data_in <= 24'b011101100100111000111011;
#10000;
	data_in <= 24'b011011000100010000110001;
#10000;
	data_in <= 24'b011001000100001100101111;
#10000;
	data_in <= 24'b010111110011111100101000;
#10000;
	data_in <= 24'b011001100100010000101101;
#10000;
	data_in <= 24'b011010100100100000110001;
#10000;
	data_in <= 24'b011001100100000100101011;
#10000;
	data_in <= 24'b011010110100011100101111;
#10000;
	data_in <= 24'b011100100100110000110100;
#10000;
	data_in <= 24'b011011000100011000101110;
#10000;
	data_in <= 24'b011000010100000100101010;
#10000;
	data_in <= 24'b011001010100011000101101;
#10000;
	data_in <= 24'b011100100101000000111000;
#10000;
	data_in <= 24'b011111110101110101000101;
#10000;
	data_in <= 24'b011011000100100000110000;
#10000;
	data_in <= 24'b011011010100101000110000;
#10000;
	data_in <= 24'b011011100100101100110001;
#10000;
	data_in <= 24'b011100010100111000110100;
#10000;
	data_in <= 24'b011000110100001100101100;
#10000;
	data_in <= 24'b011010000100100100110000;
#10000;
	data_in <= 24'b011100010101000000110110;
#10000;
	data_in <= 24'b100000100110000101000111;
#10000;
	data_in <= 24'b011100010100111000110100;
#10000;
	data_in <= 24'b011100010100111100110010;
#10000;
	data_in <= 24'b011011110100110100110000;
#10000;
	data_in <= 24'b011101010101001100110110;
#10000;
	data_in <= 24'b011011110100110100110110;
#10000;
	data_in <= 24'b011010010100011100101111;
#10000;
	data_in <= 24'b011001010100010000101010;
#10000;
	data_in <= 24'b011010100100100100101111;
#10000;
	data_in <= 24'b011010010100011100101010;
#10000;
	data_in <= 24'b011011010100101100101110;
#10000;
	data_in <= 24'b011100010100111100110010;
#10000;
	data_in <= 24'b011101010101001100110101;
#10000;
	data_in <= 24'b011011100100110000110101;
#10000;
	data_in <= 24'b011011010100101100110011;
#10000;
	data_in <= 24'b011100100101000000111000;
#10000;
	data_in <= 24'b011100000100111100110101;
#10000;
	data_in <= 24'b011101110101010000111010;
#10000;
	data_in <= 24'b011100110101000100110100;
#10000;
	data_in <= 24'b011101000101001000110101;
#10000;
	data_in <= 24'b011100100101000000110010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011001000011111100101011;
#10000;
	data_in <= 24'b011001010100000000101100;
#10000;
	data_in <= 24'b011000000011111000100111;
#10000;
	data_in <= 24'b010111110011110100100110;
#10000;
	data_in <= 24'b011000100100000000101001;
#10000;
	data_in <= 24'b011000100100001000101011;
#10000;
	data_in <= 24'b011000000100000100101000;
#10000;
	data_in <= 24'b011000010100001000101001;
#10000;
	data_in <= 24'b011011000100011000110100;
#10000;
	data_in <= 24'b011011010100100000110100;
#10000;
	data_in <= 24'b011010000100010100110001;
#10000;
	data_in <= 24'b011001010100001100101100;
#10000;
	data_in <= 24'b011000110100001100101100;
#10000;
	data_in <= 24'b011000010100000100101010;
#10000;
	data_in <= 24'b011000000100001000101001;
#10000;
	data_in <= 24'b011000100100010000101011;
#10000;
	data_in <= 24'b011010100100010100110001;
#10000;
	data_in <= 24'b011011010100100000110010;
#10000;
	data_in <= 24'b011010010100011100110000;
#10000;
	data_in <= 24'b011001100100010000101101;
#10000;
	data_in <= 24'b011000100100001000101011;
#10000;
	data_in <= 24'b011000000100000100101000;
#10000;
	data_in <= 24'b011000000100001000101001;
#10000;
	data_in <= 24'b011001000100011000101101;
#10000;
	data_in <= 24'b011010100100011000101110;
#10000;
	data_in <= 24'b011010110100011100101111;
#10000;
	data_in <= 24'b011001110100010100101101;
#10000;
	data_in <= 24'b011001100100010000101100;
#10000;
	data_in <= 24'b011001000100010100101100;
#10000;
	data_in <= 24'b011000100100001100101010;
#10000;
	data_in <= 24'b011000000100001000101001;
#10000;
	data_in <= 24'b011000100100010000101011;
#10000;
	data_in <= 24'b011100110101000000110110;
#10000;
	data_in <= 24'b011100000100110100110011;
#10000;
	data_in <= 24'b011010100100100100101111;
#10000;
	data_in <= 24'b011010100100100000110000;
#10000;
	data_in <= 24'b011010100100101100110010;
#10000;
	data_in <= 24'b011001110100011100110000;
#10000;
	data_in <= 24'b011000000100000100101010;
#10000;
	data_in <= 24'b011000010100001000101001;
#10000;
	data_in <= 24'b011101010101001100110110;
#10000;
	data_in <= 24'b011100010100111100110010;
#10000;
	data_in <= 24'b011010100100100100101111;
#10000;
	data_in <= 24'b011010110100100100110001;
#10000;
	data_in <= 24'b011011100100110000110101;
#10000;
	data_in <= 24'b011010010100100100110010;
#10000;
	data_in <= 24'b011001000100010000101101;
#10000;
	data_in <= 24'b011000110100001100101100;
#10000;
	data_in <= 24'b011100010100111100110010;
#10000;
	data_in <= 24'b011011110100110100110000;
#10000;
	data_in <= 24'b011011000100100100101111;
#10000;
	data_in <= 24'b011010110100100100110001;
#10000;
	data_in <= 24'b011011000100101000110011;
#10000;
	data_in <= 24'b011010000100011100110011;
#10000;
	data_in <= 24'b011010000100011100110011;
#10000;
	data_in <= 24'b011011000100101100110111;
#10000;
	data_in <= 24'b011100100101000000110011;
#10000;
	data_in <= 24'b011100110101000100110100;
#10000;
	data_in <= 24'b011100010100111000110100;
#10000;
	data_in <= 24'b011100000100110000110100;
#10000;
	data_in <= 24'b011011100100100100110011;
#10000;
	data_in <= 24'b011010100100011100110011;
#10000;
	data_in <= 24'b011011100100101000111000;
#10000;
	data_in <= 24'b011101110101010001000000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011000100100001100101010;
#10000;
	data_in <= 24'b011001000100010100101100;
#10000;
	data_in <= 24'b011001000100010100101100;
#10000;
	data_in <= 24'b010111110100000000100111;
#10000;
	data_in <= 24'b010111010011101100100011;
#10000;
	data_in <= 24'b010111100011110000100100;
#10000;
	data_in <= 24'b011000110011111100100111;
#10000;
	data_in <= 24'b011001010100000100101001;
#10000;
	data_in <= 24'b011001010100100000101101;
#10000;
	data_in <= 24'b011001010100100000101101;
#10000;
	data_in <= 24'b011001010100011100101100;
#10000;
	data_in <= 24'b010111110100000100100110;
#10000;
	data_in <= 24'b010111100011110100100011;
#10000;
	data_in <= 24'b010111010011110000100010;
#10000;
	data_in <= 24'b011000010011110100100101;
#10000;
	data_in <= 24'b011000100011111100100101;
#10000;
	data_in <= 24'b011001110100100100101110;
#10000;
	data_in <= 24'b011001110100100100101100;
#10000;
	data_in <= 24'b011001100100011000101001;
#10000;
	data_in <= 24'b011000100100001000100101;
#10000;
	data_in <= 24'b011000010011111100100010;
#10000;
	data_in <= 24'b011000000011111000100001;
#10000;
	data_in <= 24'b011000010011110000100010;
#10000;
	data_in <= 24'b011000010011110000100000;
#10000;
	data_in <= 24'b011001000100011000101011;
#10000;
	data_in <= 24'b011001010100010100101000;
#10000;
	data_in <= 24'b011000110100001100100110;
#10000;
	data_in <= 24'b011000010100000100100100;
#10000;
	data_in <= 24'b011000110100000100100100;
#10000;
	data_in <= 24'b011000110011111000100010;
#10000;
	data_in <= 24'b011000010011110000100000;
#10000;
	data_in <= 24'b011000010011101100011101;
#10000;
	data_in <= 24'b011000010100000000100110;
#10000;
	data_in <= 24'b011000100100000000100011;
#10000;
	data_in <= 24'b011000100100000000100010;
#10000;
	data_in <= 24'b011001000100001000100100;
#10000;
	data_in <= 24'b011010000100010000100110;
#10000;
	data_in <= 24'b011001110100001100100101;
#10000;
	data_in <= 24'b011001100100000000100010;
#10000;
	data_in <= 24'b011001000011110100011101;
#10000;
	data_in <= 24'b011000110100001000101000;
#10000;
	data_in <= 24'b011000110100000100100100;
#10000;
	data_in <= 24'b011000110100000100100100;
#10000;
	data_in <= 24'b011001100100010000100110;
#10000;
	data_in <= 24'b011010110100011100101001;
#10000;
	data_in <= 24'b011010100100011000101000;
#10000;
	data_in <= 24'b011010010100001100100011;
#10000;
	data_in <= 24'b011010000100001000100000;
#10000;
	data_in <= 24'b011010110100100100110001;
#10000;
	data_in <= 24'b011010100100100000101011;
#10000;
	data_in <= 24'b011010000100011000101001;
#10000;
	data_in <= 24'b011010100100100000101011;
#10000;
	data_in <= 24'b011011100100101000101100;
#10000;
	data_in <= 24'b011011000100100000101010;
#10000;
	data_in <= 24'b011011000100011000100110;
#10000;
	data_in <= 24'b011010110100011000100100;
#10000;
	data_in <= 24'b011100110101000100111001;
#10000;
	data_in <= 24'b011100010100111000110100;
#10000;
	data_in <= 24'b011011010100101000110000;
#10000;
	data_in <= 24'b011011010100101100101110;
#10000;
	data_in <= 24'b011011110100101100101101;
#10000;
	data_in <= 24'b011011010100101000101001;
#10000;
	data_in <= 24'b011011100100100000101000;
#10000;
	data_in <= 24'b011011010100100000100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011010010100001100101011;
#10000;
	data_in <= 24'b011001000011111000100110;
#10000;
	data_in <= 24'b011000110011110100100101;
#10000;
	data_in <= 24'b011001010011111100100111;
#10000;
	data_in <= 24'b011000110011111000100100;
#10000;
	data_in <= 24'b010111100011100100011111;
#10000;
	data_in <= 24'b010111010011100000011110;
#10000;
	data_in <= 24'b011000010011101000011110;
#10000;
	data_in <= 24'b011010000100001000101010;
#10000;
	data_in <= 24'b011001100100000100100111;
#10000;
	data_in <= 24'b011001000011111000100110;
#10000;
	data_in <= 24'b011001000011111100100101;
#10000;
	data_in <= 24'b011001100011111000100101;
#10000;
	data_in <= 24'b011000100011110100100011;
#10000;
	data_in <= 24'b011000100011101000100001;
#10000;
	data_in <= 24'b011000000011100100011101;
#10000;
	data_in <= 24'b011000110011101100100010;
#10000;
	data_in <= 24'b011001000011110100100001;
#10000;
	data_in <= 24'b011001000011110000100011;
#10000;
	data_in <= 24'b011001000011110100100001;
#10000;
	data_in <= 24'b011001110011111100100011;
#10000;
	data_in <= 24'b011010010100001000100110;
#10000;
	data_in <= 24'b011010000100000000100100;
#10000;
	data_in <= 24'b011001010011110100100000;
#10000;
	data_in <= 24'b011000000011101000011100;
#10000;
	data_in <= 24'b011000010011101100011101;
#10000;
	data_in <= 24'b011001000011110000011111;
#10000;
	data_in <= 24'b011001100011111000100001;
#10000;
	data_in <= 24'b011010000100000000100011;
#10000;
	data_in <= 24'b011010010100001000100010;
#10000;
	data_in <= 24'b011010010100001000100010;
#10000;
	data_in <= 24'b011010000100000100100001;
#10000;
	data_in <= 24'b011001010011111000011110;
#10000;
	data_in <= 24'b011001010011111000011110;
#10000;
	data_in <= 24'b011010010100000000100000;
#10000;
	data_in <= 24'b011011000100001100100011;
#10000;
	data_in <= 24'b011010110100001000100010;
#10000;
	data_in <= 24'b011001110011111000011101;
#10000;
	data_in <= 24'b011001110011111000011101;
#10000;
	data_in <= 24'b011010100100000100100000;
#10000;
	data_in <= 24'b011010010100001100100001;
#10000;
	data_in <= 24'b011001110100000100011111;
#10000;
	data_in <= 24'b011010110100001000100001;
#10000;
	data_in <= 24'b011011110100011000100101;
#10000;
	data_in <= 24'b011011100100010100100100;
#10000;
	data_in <= 24'b011010010100000100011110;
#10000;
	data_in <= 24'b011010010100000100011110;
#10000;
	data_in <= 24'b011011100100011000100011;
#10000;
	data_in <= 24'b011010110100010100100011;
#10000;
	data_in <= 24'b011010010100001100100000;
#10000;
	data_in <= 24'b011010100100010000100001;
#10000;
	data_in <= 24'b011011000100011000100011;
#10000;
	data_in <= 24'b011011100100100000100101;
#10000;
	data_in <= 24'b011011010100100000100010;
#10000;
	data_in <= 24'b011011010100100000100010;
#10000;
	data_in <= 24'b011011100100100000100101;
#10000;
	data_in <= 24'b011011100100100000100101;
#10000;
	data_in <= 24'b011011010100011100100100;
#10000;
	data_in <= 24'b011010110100010100100010;
#10000;
	data_in <= 24'b011010110100010100100010;
#10000;
	data_in <= 24'b011011100100100100100011;
#10000;
	data_in <= 24'b011100000100101100100101;
#10000;
	data_in <= 24'b011011100100100100100011;
#10000;
	data_in <= 24'b011010100100010000100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010111110011011100011010;
#10000;
	data_in <= 24'b010111110011100000011000;
#10000;
	data_in <= 24'b010111010011011000010110;
#10000;
	data_in <= 24'b010111100011011100010111;
#10000;
	data_in <= 24'b011000000011100000011011;
#10000;
	data_in <= 24'b010110110011001100010110;
#10000;
	data_in <= 24'b010110110011001100010110;
#10000;
	data_in <= 24'b011001000011111000100000;
#10000;
	data_in <= 24'b011000010011100100011100;
#10000;
	data_in <= 24'b011000110011110000011100;
#10000;
	data_in <= 24'b011000110011110000011100;
#10000;
	data_in <= 24'b011000100011101100011011;
#10000;
	data_in <= 24'b011000100011101000011101;
#10000;
	data_in <= 24'b011000000011100000011011;
#10000;
	data_in <= 24'b010111100011100000011010;
#10000;
	data_in <= 24'b011000000011101000011100;
#10000;
	data_in <= 24'b011000100011101100011011;
#10000;
	data_in <= 24'b011000110011110000011100;
#10000;
	data_in <= 24'b011001000011110000011111;
#10000;
	data_in <= 24'b011000110011101100011110;
#10000;
	data_in <= 24'b011000010011100100011100;
#10000;
	data_in <= 24'b011000110011101100011110;
#10000;
	data_in <= 24'b011000100011110000011110;
#10000;
	data_in <= 24'b010111100011100000011010;
#10000;
	data_in <= 24'b011001000011110100011101;
#10000;
	data_in <= 24'b011000100011101100011011;
#10000;
	data_in <= 24'b011000110011101100011110;
#10000;
	data_in <= 24'b011000110011101100011110;
#10000;
	data_in <= 24'b011000010011100100011100;
#10000;
	data_in <= 24'b011001010011110100100000;
#10000;
	data_in <= 24'b011001110100000100100011;
#10000;
	data_in <= 24'b011000110011110100011111;
#10000;
	data_in <= 24'b011010100100001100100011;
#10000;
	data_in <= 24'b011001010011111000011110;
#10000;
	data_in <= 24'b011001110100000000100000;
#10000;
	data_in <= 24'b011010100100001100100011;
#10000;
	data_in <= 24'b011010000100000000100011;
#10000;
	data_in <= 24'b011010100100001000100101;
#10000;
	data_in <= 24'b011011010100010100101000;
#10000;
	data_in <= 24'b011011000100010000100111;
#10000;
	data_in <= 24'b011011100100100000100110;
#10000;
	data_in <= 24'b011011000100010100100101;
#10000;
	data_in <= 24'b011011100100011100100111;
#10000;
	data_in <= 24'b011100010100101000101010;
#10000;
	data_in <= 24'b011011110100011100101010;
#10000;
	data_in <= 24'b011011010100010100101000;
#10000;
	data_in <= 24'b011011010100010100101000;
#10000;
	data_in <= 24'b011011010100010100101000;
#10000;
	data_in <= 24'b011011110100100100100111;
#10000;
	data_in <= 24'b011100100100101100101011;
#10000;
	data_in <= 24'b011100100100101100101011;
#10000;
	data_in <= 24'b011100000100100100101001;
#10000;
	data_in <= 24'b011011100100011100100111;
#10000;
	data_in <= 24'b011011000100010100100101;
#10000;
	data_in <= 24'b011010010100001000100010;
#10000;
	data_in <= 24'b011010010100001000100010;
#10000;
	data_in <= 24'b011011110100100100100111;
#10000;
	data_in <= 24'b011101110101000100101111;
#10000;
	data_in <= 24'b011100110100110000101100;
#10000;
	data_in <= 24'b011010110100010100100011;
#10000;
	data_in <= 24'b011010110100010000100100;
#10000;
	data_in <= 24'b011010110100010100100011;
#10000;
	data_in <= 24'b011010000100000100100001;
#10000;
	data_in <= 24'b011010010100001100100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011000000011100000011011;
#10000;
	data_in <= 24'b010111000011011000011000;
#10000;
	data_in <= 24'b010110100011010000010110;
#10000;
	data_in <= 24'b010110110011010000011000;
#10000;
	data_in <= 24'b010111010011011000011010;
#10000;
	data_in <= 24'b010111100011011100011011;
#10000;
	data_in <= 24'b010111010011010100011100;
#10000;
	data_in <= 24'b010110110011010000011000;
#10000;
	data_in <= 24'b011000000011101000011100;
#10000;
	data_in <= 24'b011000010011101100011101;
#10000;
	data_in <= 24'b011000110011110100011111;
#10000;
	data_in <= 24'b011001000011111000100000;
#10000;
	data_in <= 24'b011000110011110000100000;
#10000;
	data_in <= 24'b011000000011100100011101;
#10000;
	data_in <= 24'b010111010011011000011010;
#10000;
	data_in <= 24'b010110100011001100010111;
#10000;
	data_in <= 24'b010111100011100000011010;
#10000;
	data_in <= 24'b011000100011110000011110;
#10000;
	data_in <= 24'b011001010011111100100001;
#10000;
	data_in <= 24'b011001100100000000100010;
#10000;
	data_in <= 24'b011000110011110000100000;
#10000;
	data_in <= 24'b010111100011011100011011;
#10000;
	data_in <= 24'b010110110011010000011000;
#10000;
	data_in <= 24'b010110100011001100010111;
#10000;
	data_in <= 24'b011001010011111100100001;
#10000;
	data_in <= 24'b011010000100001000100100;
#10000;
	data_in <= 24'b011010100100010000100110;
#10000;
	data_in <= 24'b011010000100001000100100;
#10000;
	data_in <= 24'b011001010011111000100010;
#10000;
	data_in <= 24'b011001000011110100100001;
#10000;
	data_in <= 24'b011001000011110100100001;
#10000;
	data_in <= 24'b011001010011111000100010;
#10000;
	data_in <= 24'b011011010100011100101001;
#10000;
	data_in <= 24'b011011100100100000101010;
#10000;
	data_in <= 24'b011011000100011000101000;
#10000;
	data_in <= 24'b011010010100001100100101;
#10000;
	data_in <= 24'b011001110100000100100011;
#10000;
	data_in <= 24'b011001110100000100100011;
#10000;
	data_in <= 24'b011010010100001100100101;
#10000;
	data_in <= 24'b011010010100001100100101;
#10000;
	data_in <= 24'b011011010100011100101001;
#10000;
	data_in <= 24'b011011010100011100101001;
#10000;
	data_in <= 24'b011010110100010100100111;
#10000;
	data_in <= 24'b011001110100000100100011;
#10000;
	data_in <= 24'b011001000011111000100000;
#10000;
	data_in <= 24'b011001000011111000100000;
#10000;
	data_in <= 24'b011001000011111000100000;
#10000;
	data_in <= 24'b011000100011110000011110;
#10000;
	data_in <= 24'b011010110100010000100100;
#10000;
	data_in <= 24'b011011100100011100100111;
#10000;
	data_in <= 24'b011011010100011000100110;
#10000;
	data_in <= 24'b011010010100001000100010;
#10000;
	data_in <= 24'b011001100011111100011111;
#10000;
	data_in <= 24'b011001100011111100011111;
#10000;
	data_in <= 24'b011001010011111000011110;
#10000;
	data_in <= 24'b011000110011110000011100;
#10000;
	data_in <= 24'b011001010011111000011110;
#10000;
	data_in <= 24'b011010010100001100100001;
#10000;
	data_in <= 24'b011010100100001100100011;
#10000;
	data_in <= 24'b011001100100000000011110;
#10000;
	data_in <= 24'b011001000011110100011101;
#10000;
	data_in <= 24'b011001100100000000011110;
#10000;
	data_in <= 24'b011001110100000000100000;
#10000;
	data_in <= 24'b011001100100000000011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001011010001100100010100;
#10000;
	data_in <= 24'b001100010001110100011000;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001101110010000100011011;
#10000;
	data_in <= 24'b001110110010010100011111;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001011010001100100010100;
#10000;
	data_in <= 24'b001100000001110000010111;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001100100001111100011000;
#10000;
	data_in <= 24'b001101100010000000011010;
#10000;
	data_in <= 24'b001110100010010000011110;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001011010001100100010100;
#10000;
	data_in <= 24'b001100000001110000010111;
#10000;
	data_in <= 24'b001100010001110100011000;
#10000;
	data_in <= 24'b001100010001110100011000;
#10000;
	data_in <= 24'b001101010001111100011001;
#10000;
	data_in <= 24'b001110010010001100011101;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001011100001101000010101;
#10000;
	data_in <= 24'b001100000001110000010111;
#10000;
	data_in <= 24'b001100010001110100011000;
#10000;
	data_in <= 24'b001100100001111000011001;
#10000;
	data_in <= 24'b001101010001111100011001;
#10000;
	data_in <= 24'b001110010010001100011101;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110010010010000011100;
#10000;
	data_in <= 24'b001011110001101100010110;
#10000;
	data_in <= 24'b001100000001110000010111;
#10000;
	data_in <= 24'b001100100001111000011001;
#10000;
	data_in <= 24'b001100110001111100011010;
#10000;
	data_in <= 24'b001101100010000000011010;
#10000;
	data_in <= 24'b001110010010001100011101;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001110100010010100011101;
#10000;
	data_in <= 24'b001100000001110000010111;
#10000;
	data_in <= 24'b001100010001110100011000;
#10000;
	data_in <= 24'b001100100001111000011001;
#10000;
	data_in <= 24'b001101000010000000011011;
#10000;
	data_in <= 24'b001110000010001000011100;
#10000;
	data_in <= 24'b001110100010010000011110;
#10000;
	data_in <= 24'b001110110010011000011110;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001100010001110100011000;
#10000;
	data_in <= 24'b001100100001111000011001;
#10000;
	data_in <= 24'b001100110001111100011010;
#10000;
	data_in <= 24'b001101010010000100011100;
#10000;
	data_in <= 24'b001110010010001100011101;
#10000;
	data_in <= 24'b001110110010010100011111;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111010010100000100000;
#10000;
	data_in <= 24'b001100010001110100011000;
#10000;
	data_in <= 24'b001100100001111000011001;
#10000;
	data_in <= 24'b001100110001111100011010;
#10000;
	data_in <= 24'b001101010010000100011100;
#10000;
	data_in <= 24'b001110010010001100011101;
#10000;
	data_in <= 24'b001110110010010100011111;
#10000;
	data_in <= 24'b001111000010011100011111;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001111100010011100011111;
#10000;
	data_in <= 24'b001111110010100000100000;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000100010100100011111;
#10000;
	data_in <= 24'b010000100010100100011111;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010001100010111000100010;
#10000;
	data_in <= 24'b001111000010010100011101;
#10000;
	data_in <= 24'b001111100010011100011111;
#10000;
	data_in <= 24'b001111110010100100011110;
#10000;
	data_in <= 24'b001111110010100100011110;
#10000;
	data_in <= 24'b010000010010100000011110;
#10000;
	data_in <= 24'b010000100010100100011111;
#10000;
	data_in <= 24'b010000110010101100011111;
#10000;
	data_in <= 24'b010001110010110100100001;
#10000;
	data_in <= 24'b001111000010010100011101;
#10000;
	data_in <= 24'b001111100010011100011111;
#10000;
	data_in <= 24'b010000010010100000011110;
#10000;
	data_in <= 24'b010000100010100100011111;
#10000;
	data_in <= 24'b010000100010101000011110;
#10000;
	data_in <= 24'b010000100010101000011110;
#10000;
	data_in <= 24'b010001010010101100011111;
#10000;
	data_in <= 24'b010001110010110100100001;
#10000;
	data_in <= 24'b001111010010011000011110;
#10000;
	data_in <= 24'b001111110010100000100000;
#10000;
	data_in <= 24'b010000110010101000100000;
#10000;
	data_in <= 24'b010001000010101100100001;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010001110010110100100001;
#10000;
	data_in <= 24'b010010000010111000100010;
#10000;
	data_in <= 24'b001111110010100000100000;
#10000;
	data_in <= 24'b010000000010100100100001;
#10000;
	data_in <= 24'b010001010010110000100010;
#10000;
	data_in <= 24'b010001100010110100100011;
#10000;
	data_in <= 24'b010010000010111000100010;
#10000;
	data_in <= 24'b010010000010111000100010;
#10000;
	data_in <= 24'b010010010010111100100011;
#10000;
	data_in <= 24'b010010100011000000100100;
#10000;
	data_in <= 24'b001111110010100000100000;
#10000;
	data_in <= 24'b010000000010100100100001;
#10000;
	data_in <= 24'b010001000010101100100001;
#10000;
	data_in <= 24'b010001010010110000100010;
#10000;
	data_in <= 24'b010001110010110100100001;
#10000;
	data_in <= 24'b010010000010111000100010;
#10000;
	data_in <= 24'b010010010010111100100011;
#10000;
	data_in <= 24'b010010110011000100100101;
#10000;
	data_in <= 24'b001111110010100000100000;
#10000;
	data_in <= 24'b010000000010100100100001;
#10000;
	data_in <= 24'b010001000010101100100001;
#10000;
	data_in <= 24'b010001000010101100100001;
#10000;
	data_in <= 24'b010001100010110000100000;
#10000;
	data_in <= 24'b010001110010110100100001;
#10000;
	data_in <= 24'b010010010010111100100011;
#10000;
	data_in <= 24'b010010110011000100100101;
#10000;
	data_in <= 24'b001111110010100000100000;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010001000010101100100001;
#10000;
	data_in <= 24'b010001000010110000100000;
#10000;
	data_in <= 24'b010001100010110000100000;
#10000;
	data_in <= 24'b010001110010110100100001;
#10000;
	data_in <= 24'b010010100011000000100100;
#10000;
	data_in <= 24'b010010110011000100100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010010010010111000100000;
#10000;
	data_in <= 24'b010010010010111000100000;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010100010111100100001;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010010110011000000100010;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011000011000100100011;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010100100011011100101001;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b010100010011011000101000;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
	data_in <= 24'b010101010011100000101010;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010100000011001100100101;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010100010011010000100110;
#10000;
	data_in <= 24'b010100100011010100100111;
#10000;
	data_in <= 24'b010100110011011000101000;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010100100011010100100111;
#10000;
	data_in <= 24'b010100110011011000101000;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
	data_in <= 24'b010101100011100100101011;
#10000;
	data_in <= 24'b010110000011101100101101;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010011110011010000100110;
#10000;
	data_in <= 24'b010100100011010100100111;
#10000;
	data_in <= 24'b010100110011011000101000;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
	data_in <= 24'b010101100011100100101011;
#10000;
	data_in <= 24'b010101110011101000101100;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010100010011010000100110;
#10000;
	data_in <= 24'b010100100011010100100111;
#10000;
	data_in <= 24'b010100110011011000101000;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
	data_in <= 24'b010101010011100000101010;
#10000;
	data_in <= 24'b010101110011101000101100;
#10000;
	data_in <= 24'b010110000011101100101101;
#10000;
	data_in <= 24'b010100100011010100100111;
#10000;
	data_in <= 24'b010100110011011000101000;
#10000;
	data_in <= 24'b010101010011100000101010;
#10000;
	data_in <= 24'b010101100011100100101011;
#10000;
	data_in <= 24'b010101100011100100101011;
#10000;
	data_in <= 24'b010101110011101000101100;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010110100011110100101111;
#10000;
	data_in <= 24'b010101010011100000101010;
#10000;
	data_in <= 24'b010101100011100100101011;
#10000;
	data_in <= 24'b010101110011101000101100;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010110110011111000110000;
#10000;
	data_in <= 24'b010111000011111100110001;
#10000;
	data_in <= 24'b010111010100000000110010;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
	data_in <= 24'b010101010011100000101010;
#10000;
	data_in <= 24'b010101110011101000101100;
#10000;
	data_in <= 24'b010110000011101100101101;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010110100011110100101111;
#10000;
	data_in <= 24'b010111000011111100110001;
#10000;
	data_in <= 24'b010111010100000000110010;
#10000;
	data_in <= 24'b010100110011011000101000;
#10000;
	data_in <= 24'b010101000011011100101001;
#10000;
	data_in <= 24'b010101100011100100101011;
#10000;
	data_in <= 24'b010101110011101000101100;
#10000;
	data_in <= 24'b010110000011101100101101;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010110100011110100101111;
#10000;
	data_in <= 24'b010110100011110100101111;
#10000;
	data_in <= 24'b010101010011100000101010;
#10000;
	data_in <= 24'b010101100011100100101011;
#10000;
	data_in <= 24'b010110000011101100101101;
#10000;
	data_in <= 24'b010110010011110000101110;
#10000;
	data_in <= 24'b010110110011101100101110;
#10000;
	data_in <= 24'b010110110011101100101110;
#10000;
	data_in <= 24'b010111000011110000101111;
#10000;
	data_in <= 24'b010111010011110100110000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010110110011111000101111;
#10000;
	data_in <= 24'b010111010100000000110001;
#10000;
	data_in <= 24'b010111100100000100110010;
#10000;
	data_in <= 24'b010111110100001000110011;
#10000;
	data_in <= 24'b011000010100001000110011;
#10000;
	data_in <= 24'b011000000100000100110010;
#10000;
	data_in <= 24'b011000000100001000110001;
#10000;
	data_in <= 24'b011000000100001000110001;
#10000;
	data_in <= 24'b010110110011111000101111;
#10000;
	data_in <= 24'b010111010100000000110001;
#10000;
	data_in <= 24'b010111100100000100110010;
#10000;
	data_in <= 24'b010111110100001000110011;
#10000;
	data_in <= 24'b011000010100001000110011;
#10000;
	data_in <= 24'b011000010100001000110011;
#10000;
	data_in <= 24'b011000010100001100110010;
#10000;
	data_in <= 24'b011000010100001100110010;
#10000;
	data_in <= 24'b010111000011111100110000;
#10000;
	data_in <= 24'b010111010100000000110001;
#10000;
	data_in <= 24'b010111110100001000110011;
#10000;
	data_in <= 24'b011000000100001100110100;
#10000;
	data_in <= 24'b011000100100001100110100;
#10000;
	data_in <= 24'b011000100100001100110100;
#10000;
	data_in <= 24'b011000110100010100110100;
#10000;
	data_in <= 24'b011000110100010100110100;
#10000;
	data_in <= 24'b010111010100000000110001;
#10000;
	data_in <= 24'b010111100100000100110010;
#10000;
	data_in <= 24'b011000000100001100110100;
#10000;
	data_in <= 24'b011000010100010000110101;
#10000;
	data_in <= 24'b011000110100010000110101;
#10000;
	data_in <= 24'b011001000100010100110110;
#10000;
	data_in <= 24'b011001010100011100110110;
#10000;
	data_in <= 24'b011001100100100000110111;
#10000;
	data_in <= 24'b010111010100000000110001;
#10000;
	data_in <= 24'b010111110100001000110011;
#10000;
	data_in <= 24'b011000000100001100110100;
#10000;
	data_in <= 24'b011000010100010000110101;
#10000;
	data_in <= 24'b011001000100010100110110;
#10000;
	data_in <= 24'b011001010100011000110111;
#10000;
	data_in <= 24'b011001100100100000110111;
#10000;
	data_in <= 24'b011001110100100100111000;
#10000;
	data_in <= 24'b010111010100000000110001;
#10000;
	data_in <= 24'b010111100100000100110010;
#10000;
	data_in <= 24'b011000000100001100110100;
#10000;
	data_in <= 24'b011000010100010000110101;
#10000;
	data_in <= 24'b011000110100010000110101;
#10000;
	data_in <= 24'b011001010100011000110111;
#10000;
	data_in <= 24'b011001100100100000110111;
#10000;
	data_in <= 24'b011010000100101000111001;
#10000;
	data_in <= 24'b010111000011111100110000;
#10000;
	data_in <= 24'b010111010100000000110001;
#10000;
	data_in <= 24'b010111100100000100110010;
#10000;
	data_in <= 24'b010111110100001000110011;
#10000;
	data_in <= 24'b011000100100001100110100;
#10000;
	data_in <= 24'b011001000100010100110110;
#10000;
	data_in <= 24'b011001010100011100110110;
#10000;
	data_in <= 24'b011001110100100100111000;
#10000;
	data_in <= 24'b010111100011111100110000;
#10000;
	data_in <= 24'b010111000011111100110000;
#10000;
	data_in <= 24'b010111110100000000110001;
#10000;
	data_in <= 24'b011000000100000100110010;
#10000;
	data_in <= 24'b011000010100001000110011;
#10000;
	data_in <= 24'b011000110100010000110101;
#10000;
	data_in <= 24'b011001010100011000110111;
#10000;
	data_in <= 24'b011010000100011100111000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011000100100000100110001;
#10000;
	data_in <= 24'b011001010100010000110100;
#10000;
	data_in <= 24'b011010100100100000111000;
#10000;
	data_in <= 24'b011011010100101100111011;
#10000;
	data_in <= 24'b011011110100111000111011;
#10000;
	data_in <= 24'b011100000100111100111100;
#10000;
	data_in <= 24'b011011110100111000111011;
#10000;
	data_in <= 24'b011011110100111000111010;
#10000;
	data_in <= 24'b011001100100010100110101;
#10000;
	data_in <= 24'b011001110100011000110110;
#10000;
	data_in <= 24'b011010100100100000111000;
#10000;
	data_in <= 24'b011011010100101100111011;
#10000;
	data_in <= 24'b011100000100111100111100;
#10000;
	data_in <= 24'b011100010101000000111101;
#10000;
	data_in <= 24'b011011110100111000111011;
#10000;
	data_in <= 24'b011100000100110100111001;
#10000;
	data_in <= 24'b011001100100010100110101;
#10000;
	data_in <= 24'b011001100100010100110101;
#10000;
	data_in <= 24'b011010000100011000110110;
#10000;
	data_in <= 24'b011010100100100000111000;
#10000;
	data_in <= 24'b011011100100110100111010;
#10000;
	data_in <= 24'b011011110100111000111011;
#10000;
	data_in <= 24'b011011100100110100111010;
#10000;
	data_in <= 24'b011011100100101100110111;
#10000;
	data_in <= 24'b011001110100011000110110;
#10000;
	data_in <= 24'b011001110100011000110110;
#10000;
	data_in <= 24'b011010010100011100110111;
#10000;
	data_in <= 24'b011010110100100100111001;
#10000;
	data_in <= 24'b011011010100110000111001;
#10000;
	data_in <= 24'b011011110100111000111011;
#10000;
	data_in <= 24'b011011110100111000111011;
#10000;
	data_in <= 24'b011100000100110100111001;
#10000;
	data_in <= 24'b011011000100101100111011;
#10000;
	data_in <= 24'b011011010100110000111100;
#10000;
	data_in <= 24'b011011110100110100111101;
#10000;
	data_in <= 24'b011100000100111000111110;
#10000;
	data_in <= 24'b011100000100111100111100;
#10000;
	data_in <= 24'b011100000100111100111100;
#10000;
	data_in <= 24'b011100010101000000111101;
#10000;
	data_in <= 24'b011101000101000100111101;
#10000;
	data_in <= 24'b011011000100101100111011;
#10000;
	data_in <= 24'b011011100100110100111101;
#10000;
	data_in <= 24'b011100000100111000111110;
#10000;
	data_in <= 24'b011100000100111000111110;
#10000;
	data_in <= 24'b011011100100110100111010;
#10000;
	data_in <= 24'b011011100100110100111010;
#10000;
	data_in <= 24'b011011110100111000111011;
#10000;
	data_in <= 24'b011100110101000000111100;
#10000;
	data_in <= 24'b011010010100100000111000;
#10000;
	data_in <= 24'b011010100100100100111001;
#10000;
	data_in <= 24'b011011010100101100111011;
#10000;
	data_in <= 24'b011011010100101100111011;
#10000;
	data_in <= 24'b011011010100110000111001;
#10000;
	data_in <= 24'b011011010100110000111001;
#10000;
	data_in <= 24'b011011010100110000111001;
#10000;
	data_in <= 24'b011100000100110100111001;
#10000;
	data_in <= 24'b011010010100100000111001;
#10000;
	data_in <= 24'b011010100100100100111010;
#10000;
	data_in <= 24'b011011000100100100111011;
#10000;
	data_in <= 24'b011011100100110000111100;
#10000;
	data_in <= 24'b011100000100111000111110;
#10000;
	data_in <= 24'b011100010101000000111101;
#10000;
	data_in <= 24'b011100010100111100111111;
#10000;
	data_in <= 24'b011101010101000000111100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011110100110100110110;
#10000;
	data_in <= 24'b011100100100111000110110;
#10000;
	data_in <= 24'b011101000101000000111000;
#10000;
	data_in <= 24'b011101100101001100111001;
#10000;
	data_in <= 24'b011101010101001000111000;
#10000;
	data_in <= 24'b011100110101000100110100;
#10000;
	data_in <= 24'b011110000101001100110111;
#10000;
	data_in <= 24'b011111010101100000111100;
#10000;
	data_in <= 24'b011101010101000000111100;
#10000;
	data_in <= 24'b011101000100111100111001;
#10000;
	data_in <= 24'b011100110100111100110111;
#10000;
	data_in <= 24'b011101000101000000111000;
#10000;
	data_in <= 24'b011101100101001000111010;
#10000;
	data_in <= 24'b011101110101010000111010;
#10000;
	data_in <= 24'b011101110101001000111000;
#10000;
	data_in <= 24'b011101000100111100110101;
#10000;
	data_in <= 24'b011011110100101000110110;
#10000;
	data_in <= 24'b011100110100110000110110;
#10000;
	data_in <= 24'b011101000100110100110111;
#10000;
	data_in <= 24'b011101000100111000110110;
#10000;
	data_in <= 24'b011101100101000000111000;
#10000;
	data_in <= 24'b011101110101000100111001;
#10000;
	data_in <= 24'b011110000101001000111010;
#10000;
	data_in <= 24'b011101100101000000111000;
#10000;
	data_in <= 24'b011011110100101000110100;
#10000;
	data_in <= 24'b011100010100101000110100;
#10000;
	data_in <= 24'b011100100100101100110101;
#10000;
	data_in <= 24'b011100110100110000110110;
#10000;
	data_in <= 24'b011101010100111100110111;
#10000;
	data_in <= 24'b011101100101000000111000;
#10000;
	data_in <= 24'b011110010101001100111011;
#10000;
	data_in <= 24'b011111000101011000111110;
#10000;
	data_in <= 24'b011111110101100101000001;
#10000;
	data_in <= 24'b011110000100111100111000;
#10000;
	data_in <= 24'b011100100100100100110010;
#10000;
	data_in <= 24'b011101000100101100110100;
#10000;
	data_in <= 24'b011110000100111100111001;
#10000;
	data_in <= 24'b011110010101000000111010;
#10000;
	data_in <= 24'b011110010101000000111010;
#10000;
	data_in <= 24'b011110110101001000111100;
#10000;
	data_in <= 24'b100000010101101101000011;
#10000;
	data_in <= 24'b011110110101001100111010;
#10000;
	data_in <= 24'b011101010100110100110100;
#10000;
	data_in <= 24'b011101010100110000110101;
#10000;
	data_in <= 24'b011101100100110100110111;
#10000;
	data_in <= 24'b011101100100110100110111;
#10000;
	data_in <= 24'b011101110100111000111000;
#10000;
	data_in <= 24'b011110110101001000111100;
#10000;
	data_in <= 24'b011110000101000000110111;
#10000;
	data_in <= 24'b011110110101001100110111;
#10000;
	data_in <= 24'b011110110101001000111001;
#10000;
	data_in <= 24'b011110000100111100110110;
#10000;
	data_in <= 24'b011101110100110100110110;
#10000;
	data_in <= 24'b011110010100111100111000;
#10000;
	data_in <= 24'b011111010101001000111101;
#10000;
	data_in <= 24'b011111100101001100111110;
#10000;
	data_in <= 24'b011101110100111100110110;
#10000;
	data_in <= 24'b011111000101010000111000;
#10000;
	data_in <= 24'b011111000101001100111010;
#10000;
	data_in <= 24'b011110010100111100111000;
#10000;
	data_in <= 24'b011111000101001000111011;
#10000;
	data_in <= 24'b100001000101100101000100;
#10000;
	data_in <= 24'b100001000101100101000100;
#10000;
	data_in <= 24'b011111010101001100111100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011110010101010000111010;
#10000;
	data_in <= 24'b011110010101010000111010;
#10000;
	data_in <= 24'b011110000101001000111010;
#10000;
	data_in <= 24'b011100110100111100110111;
#10000;
	data_in <= 24'b011100010100110000110110;
#10000;
	data_in <= 24'b011100100100110100111001;
#10000;
	data_in <= 24'b011100100100110000111010;
#10000;
	data_in <= 24'b011011110100110000111000;
#10000;
	data_in <= 24'b011110010101010000111010;
#10000;
	data_in <= 24'b011110100101010100111011;
#10000;
	data_in <= 24'b011110100101010000111100;
#10000;
	data_in <= 24'b011110000101001000111010;
#10000;
	data_in <= 24'b011110000101000100111011;
#10000;
	data_in <= 24'b011101110101001000111110;
#10000;
	data_in <= 24'b011110000101000000111101;
#10000;
	data_in <= 24'b011101000100111100111011;
#10000;
	data_in <= 24'b011110110101001000111011;
#10000;
	data_in <= 24'b011111000101001100111100;
#10000;
	data_in <= 24'b011111010101010000111101;
#10000;
	data_in <= 24'b011111100101010100111110;
#10000;
	data_in <= 24'b011111110101011000111111;
#10000;
	data_in <= 24'b011111010101011001000000;
#10000;
	data_in <= 24'b011111010101010000111110;
#10000;
	data_in <= 24'b011110010101001000111100;
#10000;
	data_in <= 24'b011111000101001100111100;
#10000;
	data_in <= 24'b011111010101010000111101;
#10000;
	data_in <= 24'b011111100101010100111110;
#10000;
	data_in <= 24'b100000010101100001000001;
#10000;
	data_in <= 24'b100000110101101101000010;
#10000;
	data_in <= 24'b100000100101101001000001;
#10000;
	data_in <= 24'b011111100101010100111110;
#10000;
	data_in <= 24'b011110110101001000111011;
#10000;
	data_in <= 24'b011111110101010100111110;
#10000;
	data_in <= 24'b011111110101010100111110;
#10000;
	data_in <= 24'b100000010101100000111111;
#10000;
	data_in <= 24'b100001000101101101000010;
#10000;
	data_in <= 24'b100001010101110101000001;
#10000;
	data_in <= 24'b100000110101101100111111;
#10000;
	data_in <= 24'b011111100101011000111001;
#10000;
	data_in <= 24'b011110110101001100110111;
#10000;
	data_in <= 24'b011111100101010000111101;
#10000;
	data_in <= 24'b011111100101010100111100;
#10000;
	data_in <= 24'b100000000101011100111110;
#10000;
	data_in <= 24'b100000110101101100111111;
#10000;
	data_in <= 24'b100000110101101100111110;
#10000;
	data_in <= 24'b100000000101100100111001;
#10000;
	data_in <= 24'b011110110101010100110011;
#10000;
	data_in <= 24'b011110000101001000110000;
#10000;
	data_in <= 24'b011111010101001100111100;
#10000;
	data_in <= 24'b011111010101010000111011;
#10000;
	data_in <= 24'b100000010101011000111011;
#10000;
	data_in <= 24'b100001000101101000111101;
#10000;
	data_in <= 24'b100000110101101000111001;
#10000;
	data_in <= 24'b100000000101100000110101;
#10000;
	data_in <= 24'b011111000101010100101111;
#10000;
	data_in <= 24'b011110110101010000101110;
#10000;
	data_in <= 24'b011111100101010000111101;
#10000;
	data_in <= 24'b011111110101011100111011;
#10000;
	data_in <= 24'b100000110101100100111100;
#10000;
	data_in <= 24'b100001100101110100111101;
#10000;
	data_in <= 24'b100001110101110000111011;
#10000;
	data_in <= 24'b100001000101101000110101;
#10000;
	data_in <= 24'b100000010101100000110001;
#10000;
	data_in <= 24'b100000010101100000110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011100010100111100111000;
#10000;
	data_in <= 24'b011100110101001000111000;
#10000;
	data_in <= 24'b011100100100111100110101;
#10000;
	data_in <= 24'b011011100100110000101111;
#10000;
	data_in <= 24'b011100000100110000101110;
#10000;
	data_in <= 24'b011100010100111000101101;
#10000;
	data_in <= 24'b011100000100101000101010;
#10000;
	data_in <= 24'b011010110100011000100100;
#10000;
	data_in <= 24'b011101010101000000111010;
#10000;
	data_in <= 24'b011101010101001100111011;
#10000;
	data_in <= 24'b011101010101001000111000;
#10000;
	data_in <= 24'b011100100101000000110011;
#10000;
	data_in <= 24'b011100100100111000110000;
#10000;
	data_in <= 24'b011100100100111100101110;
#10000;
	data_in <= 24'b011101000100111000101110;
#10000;
	data_in <= 24'b011100110100111000101100;
#10000;
	data_in <= 24'b011110000101010000111100;
#10000;
	data_in <= 24'b011110010101010100111101;
#10000;
	data_in <= 24'b011110100101010100111011;
#10000;
	data_in <= 24'b011101110101001000110110;
#10000;
	data_in <= 24'b011101010100111100110001;
#10000;
	data_in <= 24'b011101000100111000101110;
#10000;
	data_in <= 24'b011101100101000000110000;
#10000;
	data_in <= 24'b011110010101010000110010;
#10000;
	data_in <= 24'b011110100101010000111100;
#10000;
	data_in <= 24'b011110100101010100111011;
#10000;
	data_in <= 24'b011110010101010000111000;
#10000;
	data_in <= 24'b011110000101001000110100;
#10000;
	data_in <= 24'b011101010100111100110001;
#10000;
	data_in <= 24'b011101000100110100101101;
#10000;
	data_in <= 24'b011101010100111100101101;
#10000;
	data_in <= 24'b011110000101001000101111;
#10000;
	data_in <= 24'b011110110101010000111000;
#10000;
	data_in <= 24'b011110010101001000110110;
#10000;
	data_in <= 24'b011101110101000100110011;
#10000;
	data_in <= 24'b011101110101000000110000;
#10000;
	data_in <= 24'b011101100101000000101110;
#10000;
	data_in <= 24'b011101100100111000101011;
#10000;
	data_in <= 24'b011101100100111100101001;
#10000;
	data_in <= 24'b011101110101000000101001;
#10000;
	data_in <= 24'b011110110101001100110110;
#10000;
	data_in <= 24'b011110010101000100110100;
#10000;
	data_in <= 24'b011110000100111100101111;
#10000;
	data_in <= 24'b011110000100111100101110;
#10000;
	data_in <= 24'b011110000101000000101101;
#10000;
	data_in <= 24'b011110110101000100101100;
#10000;
	data_in <= 24'b011110100101000100101010;
#10000;
	data_in <= 24'b011110010101000100100111;
#10000;
	data_in <= 24'b011111100101010100110100;
#10000;
	data_in <= 24'b011111010101010000110011;
#10000;
	data_in <= 24'b011111000101000100110000;
#10000;
	data_in <= 24'b011110100101000000101101;
#10000;
	data_in <= 24'b011110110101000100101100;
#10000;
	data_in <= 24'b100000000101010100101110;
#10000;
	data_in <= 24'b100000000101011000101100;
#10000;
	data_in <= 24'b011111100101010000101001;
#10000;
	data_in <= 24'b100001010101100100110100;
#10000;
	data_in <= 24'b100000110101100100110110;
#10000;
	data_in <= 24'b011111110101010100110000;
#10000;
	data_in <= 24'b011110100101000000101011;
#10000;
	data_in <= 24'b011111000101000100101010;
#10000;
	data_in <= 24'b100000000101010100101110;
#10000;
	data_in <= 24'b100000010101011100101101;
#10000;
	data_in <= 24'b011111110101010100101010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011100100100111000101010;
#10000;
	data_in <= 24'b011011110100101100100111;
#10000;
	data_in <= 24'b011011110100101100100101;
#10000;
	data_in <= 24'b011100100100111000101000;
#10000;
	data_in <= 24'b011100100100111000101000;
#10000;
	data_in <= 24'b011011110100101100100101;
#10000;
	data_in <= 24'b011011100100101000100100;
#10000;
	data_in <= 24'b011011110100101000100100;
#10000;
	data_in <= 24'b011100000100110000101000;
#10000;
	data_in <= 24'b011011010100100100100101;
#10000;
	data_in <= 24'b011011010100100100100011;
#10000;
	data_in <= 24'b011100010100110100100111;
#10000;
	data_in <= 24'b011100110100111100101001;
#10000;
	data_in <= 24'b011100010100110100100111;
#10000;
	data_in <= 24'b011100000100110000100110;
#10000;
	data_in <= 24'b011100100100110100100111;
#10000;
	data_in <= 24'b011100100100110000101001;
#10000;
	data_in <= 24'b011011110100101000100100;
#10000;
	data_in <= 24'b011011100100100100100011;
#10000;
	data_in <= 24'b011100000100101100100101;
#10000;
	data_in <= 24'b011100010100110000100110;
#10000;
	data_in <= 24'b011011110100101000100100;
#10000;
	data_in <= 24'b011011000100100000100010;
#10000;
	data_in <= 24'b011011010100100000100010;
#10000;
	data_in <= 24'b011101010101000000101010;
#10000;
	data_in <= 24'b011100100100111000100110;
#10000;
	data_in <= 24'b011100100100101100100101;
#10000;
	data_in <= 24'b011100000100110000100100;
#10000;
	data_in <= 24'b011100010100101000100100;
#10000;
	data_in <= 24'b011011000100011100100001;
#10000;
	data_in <= 24'b011010100100010100011111;
#10000;
	data_in <= 24'b011010010100010100011101;
#10000;
	data_in <= 24'b011101100100111100101000;
#10000;
	data_in <= 24'b011100110100110100100011;
#10000;
	data_in <= 24'b011100110100101000100011;
#10000;
	data_in <= 24'b011100010100101100100001;
#10000;
	data_in <= 24'b011100110100101000100011;
#10000;
	data_in <= 24'b011100000100100100100010;
#10000;
	data_in <= 24'b011011100100011100100000;
#10000;
	data_in <= 24'b011011100100011100100000;
#10000;
	data_in <= 24'b011110000100111000100100;
#10000;
	data_in <= 24'b011101000100110100100001;
#10000;
	data_in <= 24'b011101000100101000100000;
#10000;
	data_in <= 24'b011100100100101000100000;
#10000;
	data_in <= 24'b011101000100101000100000;
#10000;
	data_in <= 24'b011100100100101000100000;
#10000;
	data_in <= 24'b011100010100100100011111;
#10000;
	data_in <= 24'b011100000100100000011110;
#10000;
	data_in <= 24'b011110100100111100100100;
#10000;
	data_in <= 24'b011110000100111100100010;
#10000;
	data_in <= 24'b011101100100101100100000;
#10000;
	data_in <= 24'b011101000100101000011111;
#10000;
	data_in <= 24'b011101010100101000011111;
#10000;
	data_in <= 24'b011101000100101000011111;
#10000;
	data_in <= 24'b011100110100100100011110;
#10000;
	data_in <= 24'b011100010100011100011100;
#10000;
	data_in <= 24'b011111000101000100100110;
#10000;
	data_in <= 24'b011110100100111100100100;
#10000;
	data_in <= 24'b011110000100110100100010;
#10000;
	data_in <= 24'b011101110100110000100001;
#10000;
	data_in <= 24'b011110000100110100100010;
#10000;
	data_in <= 24'b011110010100111000100011;
#10000;
	data_in <= 24'b011101110100110100100010;
#10000;
	data_in <= 24'b011101100100110100100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011101010100111100101100;
#10000;
	data_in <= 24'b011101000100110000101001;
#10000;
	data_in <= 24'b011101000100101100101010;
#10000;
	data_in <= 24'b011100010100100100100110;
#10000;
	data_in <= 24'b011010110100001000100001;
#10000;
	data_in <= 24'b011010000100000000011101;
#10000;
	data_in <= 24'b011010100100000100100000;
#10000;
	data_in <= 24'b011011000100010000100001;
#10000;
	data_in <= 24'b100001100101111100111001;
#10000;
	data_in <= 24'b011110000101000100101011;
#10000;
	data_in <= 24'b011011010100010100100010;
#10000;
	data_in <= 24'b011010010100001000011100;
#10000;
	data_in <= 24'b011010110100001100100000;
#10000;
	data_in <= 24'b011011100100011100100001;
#10000;
	data_in <= 24'b011011100100011000100011;
#10000;
	data_in <= 24'b011010100100001100011101;
#10000;
	data_in <= 24'b011110100101001100101101;
#10000;
	data_in <= 24'b011100110100101000100011;
#10000;
	data_in <= 24'b011011000100001000011101;
#10000;
	data_in <= 24'b011011000100001100011100;
#10000;
	data_in <= 24'b011011000100001000011101;
#10000;
	data_in <= 24'b011011110100011000011111;
#10000;
	data_in <= 24'b011011110100010100100000;
#10000;
	data_in <= 24'b011011000100001100011100;
#10000;
	data_in <= 24'b011010110100001000011011;
#10000;
	data_in <= 24'b011010110100001100011001;
#10000;
	data_in <= 24'b011011100100010100011110;
#10000;
	data_in <= 24'b011100000100100000011110;
#10000;
	data_in <= 24'b011011000100010000011010;
#10000;
	data_in <= 24'b011010110100001100011001;
#10000;
	data_in <= 24'b011011010100010100011011;
#10000;
	data_in <= 24'b011100000100011000011100;
#10000;
	data_in <= 24'b011100010100100100011111;
#10000;
	data_in <= 24'b011011110100010100011010;
#10000;
	data_in <= 24'b011011110100010100011011;
#10000;
	data_in <= 24'b011100000100011000011011;
#10000;
	data_in <= 24'b011011100100010000011001;
#10000;
	data_in <= 24'b011011100100010000011001;
#10000;
	data_in <= 24'b011011110100010100011010;
#10000;
	data_in <= 24'b011011110100010000011001;
#10000;
	data_in <= 24'b011101000100101000011111;
#10000;
	data_in <= 24'b011011110100011000011001;
#10000;
	data_in <= 24'b011011100100010000011001;
#10000;
	data_in <= 24'b011011110100011000011001;
#10000;
	data_in <= 24'b011011100100010100011000;
#10000;
	data_in <= 24'b011011100100010100011000;
#10000;
	data_in <= 24'b011011110100010100011000;
#10000;
	data_in <= 24'b011011010100001100010110;
#10000;
	data_in <= 24'b011011110100011000011001;
#10000;
	data_in <= 24'b011011110100010100010110;
#10000;
	data_in <= 24'b011100010100011100011010;
#10000;
	data_in <= 24'b011100100100100000011001;
#10000;
	data_in <= 24'b011011110100010100010110;
#10000;
	data_in <= 24'b011011010100001100010100;
#10000;
	data_in <= 24'b011011100100010000010101;
#10000;
	data_in <= 24'b011011010100001100010100;
#10000;
	data_in <= 24'b011110010100111100100010;
#10000;
	data_in <= 24'b011101000100101000011011;
#10000;
	data_in <= 24'b011100110100100100011010;
#10000;
	data_in <= 24'b011100110100100100011010;
#10000;
	data_in <= 24'b011100010100011100011000;
#10000;
	data_in <= 24'b011100010100011100011000;
#10000;
	data_in <= 24'b011100010100011100011000;
#10000;
	data_in <= 24'b011011110100010100010110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011000100001100100010;
#10000;
	data_in <= 24'b011011000100010000100001;
#10000;
	data_in <= 24'b011010110100001000100001;
#10000;
	data_in <= 24'b011010110100001100100000;
#10000;
	data_in <= 24'b011011000100001100100010;
#10000;
	data_in <= 24'b011011000100010000100001;
#10000;
	data_in <= 24'b011010100100000100100000;
#10000;
	data_in <= 24'b011001100011111000011011;
#10000;
	data_in <= 24'b011011010100011000100000;
#10000;
	data_in <= 24'b011011010100011000100000;
#10000;
	data_in <= 24'b011011100100010000011111;
#10000;
	data_in <= 24'b011010110100010000011110;
#10000;
	data_in <= 24'b011011000100001000011101;
#10000;
	data_in <= 24'b011010100100001100011101;
#10000;
	data_in <= 24'b011010100100000000011011;
#10000;
	data_in <= 24'b011001000011110100010111;
#10000;
	data_in <= 24'b011010110100001000011011;
#10000;
	data_in <= 24'b011011000100001100011100;
#10000;
	data_in <= 24'b011011100100001100011100;
#10000;
	data_in <= 24'b011010100100000100011010;
#10000;
	data_in <= 24'b011010110100000000011001;
#10000;
	data_in <= 24'b011010000011111100011000;
#10000;
	data_in <= 24'b011010000011110100010110;
#10000;
	data_in <= 24'b011001000011101100010100;
#10000;
	data_in <= 24'b011010010011111100010101;
#10000;
	data_in <= 24'b011010100100000000010101;
#10000;
	data_in <= 24'b011010110100000100010111;
#10000;
	data_in <= 24'b011010100100000000010101;
#10000;
	data_in <= 24'b011010010011111100010101;
#10000;
	data_in <= 24'b011010000011111000010011;
#10000;
	data_in <= 24'b011001110011110100010011;
#10000;
	data_in <= 24'b011001100011110000010001;
#10000;
	data_in <= 24'b011010110100000000010101;
#10000;
	data_in <= 24'b011010110100000100010100;
#10000;
	data_in <= 24'b011011000100000100010110;
#10000;
	data_in <= 24'b011011000100001000010101;
#10000;
	data_in <= 24'b011010110100000000010101;
#10000;
	data_in <= 24'b011010100100000000010011;
#10000;
	data_in <= 24'b011010010011111000010011;
#10000;
	data_in <= 24'b011010010011111100010010;
#10000;
	data_in <= 24'b011011100100010000010111;
#10000;
	data_in <= 24'b011011010100001100010100;
#10000;
	data_in <= 24'b011011000100001000010101;
#10000;
	data_in <= 24'b011011000100001000010011;
#10000;
	data_in <= 24'b011010110100000100010100;
#10000;
	data_in <= 24'b011010010011111100010000;
#10000;
	data_in <= 24'b011010000011111000010001;
#10000;
	data_in <= 24'b011010000011111000001111;
#10000;
	data_in <= 24'b011100100100011000010111;
#10000;
	data_in <= 24'b011011110100010000010011;
#10000;
	data_in <= 24'b011011100100001000010011;
#10000;
	data_in <= 24'b011011100100001100010010;
#10000;
	data_in <= 24'b011011010100000100010010;
#10000;
	data_in <= 24'b011010110100000000001111;
#10000;
	data_in <= 24'b011010010011110100001110;
#10000;
	data_in <= 24'b011010000011110100001100;
#10000;
	data_in <= 24'b011101000100100000011001;
#10000;
	data_in <= 24'b011100000100010100010100;
#10000;
	data_in <= 24'b011011100100001000010011;
#10000;
	data_in <= 24'b011011110100010000010011;
#10000;
	data_in <= 24'b011011110100010000010011;
#10000;
	data_in <= 24'b011011010100001000010001;
#10000;
	data_in <= 24'b011010110100000000001111;
#10000;
	data_in <= 24'b011010100011111100001110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001100010001111000011001;
#10000;
	data_in <= 24'b001100100001111100011010;
#10000;
	data_in <= 24'b001101000010000100011100;
#10000;
	data_in <= 24'b001101100010001100011110;
#10000;
	data_in <= 24'b001110010010011000011111;
#10000;
	data_in <= 24'b001110100010011100100000;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b001100010001111000011001;
#10000;
	data_in <= 24'b001100100001111100011010;
#10000;
	data_in <= 24'b001101010010001000011101;
#10000;
	data_in <= 24'b001101100010001100011110;
#10000;
	data_in <= 24'b001110010010011000011111;
#10000;
	data_in <= 24'b001110100010011100100000;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b001100010001111000011001;
#10000;
	data_in <= 24'b001100110010000000011011;
#10000;
	data_in <= 24'b001101010010001000011101;
#10000;
	data_in <= 24'b001101110010010000011111;
#10000;
	data_in <= 24'b001110010010011000011111;
#10000;
	data_in <= 24'b001110110010100000100001;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b001100010001111000011001;
#10000;
	data_in <= 24'b001100110010000000011011;
#10000;
	data_in <= 24'b001101010010001000011101;
#10000;
	data_in <= 24'b001101110010010000011111;
#10000;
	data_in <= 24'b001110010010011000011111;
#10000;
	data_in <= 24'b001110110010100000100001;
#10000;
	data_in <= 24'b001111100010100100100001;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b001100000001110100011000;
#10000;
	data_in <= 24'b001100100001111100011010;
#10000;
	data_in <= 24'b001101000010000100011100;
#10000;
	data_in <= 24'b001101100010001100011110;
#10000;
	data_in <= 24'b001110000010010100011110;
#10000;
	data_in <= 24'b001110100010011100100000;
#10000;
	data_in <= 24'b001111100010100000100010;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b001011110001110000010111;
#10000;
	data_in <= 24'b001100010001111000011001;
#10000;
	data_in <= 24'b001100110010000000011011;
#10000;
	data_in <= 24'b001101010010001000011101;
#10000;
	data_in <= 24'b001101110010010000011101;
#10000;
	data_in <= 24'b001110010010011000011111;
#10000;
	data_in <= 24'b001111000010011000100000;
#10000;
	data_in <= 24'b001111100010100000100010;
#10000;
	data_in <= 24'b001011100001101100010110;
#10000;
	data_in <= 24'b001011110001110000010111;
#10000;
	data_in <= 24'b001100100001111100011010;
#10000;
	data_in <= 24'b001100110010000000011011;
#10000;
	data_in <= 24'b001101100010001000011101;
#10000;
	data_in <= 24'b001101110010001100011110;
#10000;
	data_in <= 24'b001110010010011000011111;
#10000;
	data_in <= 24'b001110100010011100100000;
#10000;
	data_in <= 24'b001011010001101000010101;
#10000;
	data_in <= 24'b001011110001110000010111;
#10000;
	data_in <= 24'b001100010001111000011001;
#10000;
	data_in <= 24'b001100110010000000011011;
#10000;
	data_in <= 24'b001101010010000100011100;
#10000;
	data_in <= 24'b001101110010001100011110;
#10000;
	data_in <= 24'b001110000010010100011110;
#10000;
	data_in <= 24'b001110010010011000011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001111100010100000011101;
#10000;
	data_in <= 24'b010000000010101000011111;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b010001110010111100100011;
#10000;
	data_in <= 24'b010001110011000000100001;
#10000;
	data_in <= 24'b010010110011000100100011;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010000110010110100100001;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b010001110010111100100011;
#10000;
	data_in <= 24'b010010000011000100100010;
#10000;
	data_in <= 24'b010011000011001000100100;
#10000;
	data_in <= 24'b010011010011001100100101;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010001000010111000100010;
#10000;
	data_in <= 24'b010001110010111100100011;
#10000;
	data_in <= 24'b010010000011000000100100;
#10000;
	data_in <= 24'b010010010011000100100101;
#10000;
	data_in <= 24'b010011000011001000100110;
#10000;
	data_in <= 24'b010001010010111000100110;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010000110010110100100010;
#10000;
	data_in <= 24'b010001110010111100100011;
#10000;
	data_in <= 24'b010010000011000000100100;
#10000;
	data_in <= 24'b010010010011000100100101;
#10000;
	data_in <= 24'b010010010011000100100101;
#10000;
	data_in <= 24'b010000010010110000100100;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b010000100010110000100001;
#10000;
	data_in <= 24'b010001000010111000100011;
#10000;
	data_in <= 24'b010001100011000000100101;
#10000;
	data_in <= 24'b010001110011000100100110;
#10000;
	data_in <= 24'b010010010011000100100101;
#10000;
	data_in <= 24'b010010000011000000100100;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000110010110000100100;
#10000;
	data_in <= 24'b010001010010111100100100;
#10000;
	data_in <= 24'b010001100011000000100101;
#10000;
	data_in <= 24'b010010000011001000100111;
#10000;
	data_in <= 24'b010010100011000100100111;
#10000;
	data_in <= 24'b010010100011001000100110;
#10000;
	data_in <= 24'b001111100010100000100010;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b010000100010110100100101;
#10000;
	data_in <= 24'b010000110010111000100110;
#10000;
	data_in <= 24'b010001000011000000100101;
#10000;
	data_in <= 24'b010010000011001000100111;
#10000;
	data_in <= 24'b010010010011001100101000;
#10000;
	data_in <= 24'b001111000010100100100010;
#10000;
	data_in <= 24'b001111100010100000100010;
#10000;
	data_in <= 24'b001111110010101000100010;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b010000000010101100100011;
#10000;
	data_in <= 24'b010000100010110100100101;
#10000;
	data_in <= 24'b010001010011000000101000;
#10000;
	data_in <= 24'b010010010011001100101000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100100011010000101001;
#10000;
	data_in <= 24'b010100010011001100101000;
#10000;
	data_in <= 24'b010100110011001100101000;
#10000;
	data_in <= 24'b010100010011001100101000;
#10000;
	data_in <= 24'b010100110011001100101000;
#10000;
	data_in <= 24'b010101010011010100101010;
#10000;
	data_in <= 24'b010101100011011000101011;
#10000;
	data_in <= 24'b010101110011011100101100;
#10000;
	data_in <= 24'b010100010011001100101000;
#10000;
	data_in <= 24'b010100010011001100101000;
#10000;
	data_in <= 24'b010101000011010000101001;
#10000;
	data_in <= 24'b010100100011010000101001;
#10000;
	data_in <= 24'b010101010011010100101010;
#10000;
	data_in <= 24'b010101000011011000101011;
#10000;
	data_in <= 24'b010101110011011100101100;
#10000;
	data_in <= 24'b010101100011100000101101;
#10000;
	data_in <= 24'b010011010011001000100100;
#10000;
	data_in <= 24'b010011100011001100100101;
#10000;
	data_in <= 24'b010100100011010000101001;
#10000;
	data_in <= 24'b010100010011010100101010;
#10000;
	data_in <= 24'b010101000011011000101011;
#10000;
	data_in <= 24'b010100110011011100101100;
#10000;
	data_in <= 24'b010101010011011100101100;
#10000;
	data_in <= 24'b010101000011100000101101;
#10000;
	data_in <= 24'b010010110011000100100011;
#10000;
	data_in <= 24'b010011000011001000100100;
#10000;
	data_in <= 24'b010011100011001000100111;
#10000;
	data_in <= 24'b010011110011010100101001;
#10000;
	data_in <= 24'b010100010011010100101010;
#10000;
	data_in <= 24'b010100010011011100101011;
#10000;
	data_in <= 24'b010100110011011100101100;
#10000;
	data_in <= 24'b010100100011100000101100;
#10000;
	data_in <= 24'b010010100011001000100110;
#10000;
	data_in <= 24'b010010100011001000100110;
#10000;
	data_in <= 24'b010011010011001100100111;
#10000;
	data_in <= 24'b010011000011010000101000;
#10000;
	data_in <= 24'b010011110011010000101010;
#10000;
	data_in <= 24'b010011110011011000101100;
#10000;
	data_in <= 24'b010100100011011100101101;
#10000;
	data_in <= 24'b010100010011100000101110;
#10000;
	data_in <= 24'b010011000011010000101000;
#10000;
	data_in <= 24'b010011000011010000101000;
#10000;
	data_in <= 24'b010011000011010000101000;
#10000;
	data_in <= 24'b010011010011010100101001;
#10000;
	data_in <= 24'b010011100011010100101011;
#10000;
	data_in <= 24'b010100000011011100101101;
#10000;
	data_in <= 24'b010100010011100000101110;
#10000;
	data_in <= 24'b010100100011100100101111;
#10000;
	data_in <= 24'b010010110011010100101001;
#10000;
	data_in <= 24'b010010110011010100101001;
#10000;
	data_in <= 24'b010011000011011000101011;
#10000;
	data_in <= 24'b010011010011011100101100;
#10000;
	data_in <= 24'b010011100011011100101111;
#10000;
	data_in <= 24'b010011110011100000110000;
#10000;
	data_in <= 24'b010011110011100000110000;
#10000;
	data_in <= 24'b010011110011100000110000;
#10000;
	data_in <= 24'b010010100011010000101001;
#10000;
	data_in <= 24'b010010110011010100101001;
#10000;
	data_in <= 24'b010011010011011100101100;
#10000;
	data_in <= 24'b010011100011100000101101;
#10000;
	data_in <= 24'b010011110011100000110000;
#10000;
	data_in <= 24'b010011110011100000110000;
#10000;
	data_in <= 24'b010011100011011100101111;
#10000;
	data_in <= 24'b010011100011011100101111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010110010011100100101110;
#10000;
	data_in <= 24'b010110010011100100101110;
#10000;
	data_in <= 24'b010110010011100100101100;
#10000;
	data_in <= 24'b010110100011101000101101;
#10000;
	data_in <= 24'b010111010011110000101101;
#10000;
	data_in <= 24'b010111100011110100101110;
#10000;
	data_in <= 24'b010111110011111000101111;
#10000;
	data_in <= 24'b011000000011111100110000;
#10000;
	data_in <= 24'b010110010011100100101110;
#10000;
	data_in <= 24'b010110010011100100101110;
#10000;
	data_in <= 24'b010110100011101000101101;
#10000;
	data_in <= 24'b010111000011101000101101;
#10000;
	data_in <= 24'b010111010011101100101110;
#10000;
	data_in <= 24'b010111110011111000101111;
#10000;
	data_in <= 24'b011000000011111100110000;
#10000;
	data_in <= 24'b011000000011111100110000;
#10000;
	data_in <= 24'b010110000011101000101111;
#10000;
	data_in <= 24'b010110000011101000101111;
#10000;
	data_in <= 24'b010110000011101000101111;
#10000;
	data_in <= 24'b010110110011101100101110;
#10000;
	data_in <= 24'b010111000011110000101111;
#10000;
	data_in <= 24'b010111010011110100110000;
#10000;
	data_in <= 24'b010111100011111000110001;
#10000;
	data_in <= 24'b010111100011111000110001;
#10000;
	data_in <= 24'b010101100011101000101111;
#10000;
	data_in <= 24'b010101100011101000101111;
#10000;
	data_in <= 24'b010101100011101000101111;
#10000;
	data_in <= 24'b010110010011101100110000;
#10000;
	data_in <= 24'b010110100011110000110001;
#10000;
	data_in <= 24'b010110100011110100101111;
#10000;
	data_in <= 24'b010111010011110100110000;
#10000;
	data_in <= 24'b010111100011111000110001;
#10000;
	data_in <= 24'b010101010011101000110000;
#10000;
	data_in <= 24'b010101010011101000110000;
#10000;
	data_in <= 24'b010101010011101000110000;
#10000;
	data_in <= 24'b010101100011100100110000;
#10000;
	data_in <= 24'b010101110011101000110001;
#10000;
	data_in <= 24'b010110000011110000110001;
#10000;
	data_in <= 24'b010110110011110100110010;
#10000;
	data_in <= 24'b010110110011111000110000;
#10000;
	data_in <= 24'b010100100011100100101111;
#10000;
	data_in <= 24'b010100100011100100101111;
#10000;
	data_in <= 24'b010101010011100100110010;
#10000;
	data_in <= 24'b010101010011101000110000;
#10000;
	data_in <= 24'b010101100011100100110000;
#10000;
	data_in <= 24'b010101110011101000110001;
#10000;
	data_in <= 24'b010101110011101000110001;
#10000;
	data_in <= 24'b010110000011110000110001;
#10000;
	data_in <= 24'b010100000011100100110001;
#10000;
	data_in <= 24'b010100000011100100110001;
#10000;
	data_in <= 24'b010100100011100000110010;
#10000;
	data_in <= 24'b010100100011100000110001;
#10000;
	data_in <= 24'b010101000011100000110001;
#10000;
	data_in <= 24'b010101010011100100110010;
#10000;
	data_in <= 24'b010101100011100100110010;
#10000;
	data_in <= 24'b010101110011101000110001;
#10000;
	data_in <= 24'b010011110011011100110001;
#10000;
	data_in <= 24'b010011110011011100110001;
#10000;
	data_in <= 24'b010100010011011100110001;
#10000;
	data_in <= 24'b010100010011011100110001;
#10000;
	data_in <= 24'b010101000011011100110010;
#10000;
	data_in <= 24'b010101000011100000110001;
#10000;
	data_in <= 24'b010101100011100100110010;
#10000;
	data_in <= 24'b010101100011100100110010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011000010100000000110001;
#10000;
	data_in <= 24'b011000000100000100110010;
#10000;
	data_in <= 24'b011000100100000100110010;
#10000;
	data_in <= 24'b011000110100001000110011;
#10000;
	data_in <= 24'b011001000100001000110101;
#10000;
	data_in <= 24'b011001010100001100110110;
#10000;
	data_in <= 24'b011001110100010100111000;
#10000;
	data_in <= 24'b011010100100011100111010;
#10000;
	data_in <= 24'b011000100100000100110010;
#10000;
	data_in <= 24'b011000110100001000110011;
#10000;
	data_in <= 24'b011000110100001000110011;
#10000;
	data_in <= 24'b011001000100001100110100;
#10000;
	data_in <= 24'b011001010100001100110110;
#10000;
	data_in <= 24'b011001100100010000110111;
#10000;
	data_in <= 24'b011010010100010100111011;
#10000;
	data_in <= 24'b011010110100011100111101;
#10000;
	data_in <= 24'b011000000100000100110010;
#10000;
	data_in <= 24'b011000010100001000110011;
#10000;
	data_in <= 24'b011001000100001000110101;
#10000;
	data_in <= 24'b011001010100001100110110;
#10000;
	data_in <= 24'b011001010100001100110110;
#10000;
	data_in <= 24'b011001110100010100111000;
#10000;
	data_in <= 24'b011010100100011000111100;
#10000;
	data_in <= 24'b011010110100011100111101;
#10000;
	data_in <= 24'b010111110011111100110010;
#10000;
	data_in <= 24'b011000000100000100110010;
#10000;
	data_in <= 24'b011000110100000100110100;
#10000;
	data_in <= 24'b011001000100001000110101;
#10000;
	data_in <= 24'b011001010100001100110110;
#10000;
	data_in <= 24'b011001100100010000110111;
#10000;
	data_in <= 24'b011010010100010100111011;
#10000;
	data_in <= 24'b011010100100011000111100;
#10000;
	data_in <= 24'b010111000011111100110001;
#10000;
	data_in <= 24'b010111010100000000110010;
#10000;
	data_in <= 24'b011000000100000000110101;
#10000;
	data_in <= 24'b011000010100000100110110;
#10000;
	data_in <= 24'b011000100100001000110111;
#10000;
	data_in <= 24'b011001000100010000111001;
#10000;
	data_in <= 24'b011001110100010000111010;
#10000;
	data_in <= 24'b011010010100011000111100;
#10000;
	data_in <= 24'b010110110011110100110010;
#10000;
	data_in <= 24'b010111000011111000110011;
#10000;
	data_in <= 24'b010111100100000000110101;
#10000;
	data_in <= 24'b011000010100000100110110;
#10000;
	data_in <= 24'b011000100100001000110111;
#10000;
	data_in <= 24'b011000110100001100111000;
#10000;
	data_in <= 24'b011001110100010000111010;
#10000;
	data_in <= 24'b011010000100010100111011;
#10000;
	data_in <= 24'b010110000011101100110010;
#10000;
	data_in <= 24'b010110010011110000110011;
#10000;
	data_in <= 24'b010110100011110100110100;
#10000;
	data_in <= 24'b010111100011111100110110;
#10000;
	data_in <= 24'b011000010100000000110111;
#10000;
	data_in <= 24'b011000100100000100111000;
#10000;
	data_in <= 24'b011001100100001000111010;
#10000;
	data_in <= 24'b011001110100001100111011;
#10000;
	data_in <= 24'b010101100011100100110010;
#10000;
	data_in <= 24'b010101110011101000110001;
#10000;
	data_in <= 24'b010110010011110000110011;
#10000;
	data_in <= 24'b010110100011110100110100;
#10000;
	data_in <= 24'b010111010011111000110101;
#10000;
	data_in <= 24'b011000010100000000110111;
#10000;
	data_in <= 24'b011001000100000000111000;
#10000;
	data_in <= 24'b011001010100000100111001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011010110100100000111011;
#10000;
	data_in <= 24'b011010110100100000111011;
#10000;
	data_in <= 24'b011011010100011100111011;
#10000;
	data_in <= 24'b011011110100101000111100;
#10000;
	data_in <= 24'b011100100100110100111111;
#10000;
	data_in <= 24'b011101000101000001000000;
#10000;
	data_in <= 24'b011101000100111101000001;
#10000;
	data_in <= 24'b011101100101000000111110;
#10000;
	data_in <= 24'b011011000100100000111110;
#10000;
	data_in <= 24'b011011000100100000111110;
#10000;
	data_in <= 24'b011011100100100000111100;
#10000;
	data_in <= 24'b011100000100101000111110;
#10000;
	data_in <= 24'b011100100100110100111111;
#10000;
	data_in <= 24'b011101000100111101000001;
#10000;
	data_in <= 24'b011101110101000001000010;
#10000;
	data_in <= 24'b011101110101000001000001;
#10000;
	data_in <= 24'b011011000100100000111110;
#10000;
	data_in <= 24'b011011000100100000111110;
#10000;
	data_in <= 24'b011011110100100100111101;
#10000;
	data_in <= 24'b011100010100101100111111;
#10000;
	data_in <= 24'b011101010100111001000000;
#10000;
	data_in <= 24'b011101100100111101000001;
#10000;
	data_in <= 24'b011101110101000001000010;
#10000;
	data_in <= 24'b011101110101000001000001;
#10000;
	data_in <= 24'b011011000100100000111110;
#10000;
	data_in <= 24'b011011010100100100111111;
#10000;
	data_in <= 24'b011100000100101000111110;
#10000;
	data_in <= 24'b011100010100101100111111;
#10000;
	data_in <= 24'b011101010100111001000000;
#10000;
	data_in <= 24'b011101100100111101000001;
#10000;
	data_in <= 24'b011101110101000001000010;
#10000;
	data_in <= 24'b011101110101000001000001;
#10000;
	data_in <= 24'b011010110100011100111101;
#10000;
	data_in <= 24'b011011000100100000111110;
#10000;
	data_in <= 24'b011100000100101000111110;
#10000;
	data_in <= 24'b011100010100101100111111;
#10000;
	data_in <= 24'b011101010100111001000000;
#10000;
	data_in <= 24'b011101100100111101000001;
#10000;
	data_in <= 24'b011101110101000001000010;
#10000;
	data_in <= 24'b011101110101000001000010;
#10000;
	data_in <= 24'b011010100100011000111100;
#10000;
	data_in <= 24'b011010110100011100111101;
#10000;
	data_in <= 24'b011011110100100100111101;
#10000;
	data_in <= 24'b011100010100101100111111;
#10000;
	data_in <= 24'b011101000100110001000000;
#10000;
	data_in <= 24'b011101010100111001000000;
#10000;
	data_in <= 24'b011101100100111101000001;
#10000;
	data_in <= 24'b011101110101000001000010;
#10000;
	data_in <= 24'b011010000100010000111010;
#10000;
	data_in <= 24'b011010100100011000111100;
#10000;
	data_in <= 24'b011011100100011100111110;
#10000;
	data_in <= 24'b011100000100100101000000;
#10000;
	data_in <= 24'b011100010100101001000001;
#10000;
	data_in <= 24'b011100100100110001000000;
#10000;
	data_in <= 24'b011101000100111001000010;
#10000;
	data_in <= 24'b011101000100111001000010;
#10000;
	data_in <= 24'b011001110100001000111010;
#10000;
	data_in <= 24'b011010010100010100111011;
#10000;
	data_in <= 24'b011010110100011000111110;
#10000;
	data_in <= 24'b011011010100100100111111;
#10000;
	data_in <= 24'b011100010100101001000010;
#10000;
	data_in <= 24'b011100000100110001000010;
#10000;
	data_in <= 24'b011100110100110001000011;
#10000;
	data_in <= 24'b011101000100110101000100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011110110101001000111100;
#10000;
	data_in <= 24'b011111000101001100111100;
#10000;
	data_in <= 24'b011110110101001000111100;
#10000;
	data_in <= 24'b011110110101001000111100;
#10000;
	data_in <= 24'b011111010101010000111110;
#10000;
	data_in <= 24'b100000000101011101000001;
#10000;
	data_in <= 24'b100000100101100101000011;
#10000;
	data_in <= 24'b100000100101100101000010;
#10000;
	data_in <= 24'b011111000101001000111111;
#10000;
	data_in <= 24'b011111100101010100111111;
#10000;
	data_in <= 24'b011111110101010101000010;
#10000;
	data_in <= 24'b011111110101010101000010;
#10000;
	data_in <= 24'b011111110101011101000100;
#10000;
	data_in <= 24'b100000110101101101001000;
#10000;
	data_in <= 24'b100010000101111101001001;
#10000;
	data_in <= 24'b100010000101111101001000;
#10000;
	data_in <= 24'b011111000101000101000000;
#10000;
	data_in <= 24'b011111110101010101000010;
#10000;
	data_in <= 24'b100000010101011101000100;
#10000;
	data_in <= 24'b100000100101100001000101;
#10000;
	data_in <= 24'b100000010101100101000110;
#10000;
	data_in <= 24'b100001000101110001001001;
#10000;
	data_in <= 24'b100010010110000001001010;
#10000;
	data_in <= 24'b100010100110000101001010;
#10000;
	data_in <= 24'b011110100101001001000000;
#10000;
	data_in <= 24'b011111110101010101000010;
#10000;
	data_in <= 24'b100000010101011101000100;
#10000;
	data_in <= 24'b100000100101100001000101;
#10000;
	data_in <= 24'b100000000101100001000101;
#10000;
	data_in <= 24'b100000100101101001000111;
#10000;
	data_in <= 24'b100001100101110101000111;
#10000;
	data_in <= 24'b100001100101110101000110;
#10000;
	data_in <= 24'b011110100101000101000010;
#10000;
	data_in <= 24'b011111010101010101000011;
#10000;
	data_in <= 24'b011111110101011101000101;
#10000;
	data_in <= 24'b100000000101100001000110;
#10000;
	data_in <= 24'b100000000101100001000110;
#10000;
	data_in <= 24'b100000010101100101000110;
#10000;
	data_in <= 24'b100001000101101101000101;
#10000;
	data_in <= 24'b100001000101101101000100;
#10000;
	data_in <= 24'b011110010100111101000010;
#10000;
	data_in <= 24'b011110110101001001000011;
#10000;
	data_in <= 24'b011111000101001101000100;
#10000;
	data_in <= 24'b011111010101010101000011;
#10000;
	data_in <= 24'b011111110101011101000101;
#10000;
	data_in <= 24'b100000010101100101000110;
#10000;
	data_in <= 24'b100001000101101001000111;
#10000;
	data_in <= 24'b100000110101101001000011;
#10000;
	data_in <= 24'b011101100100111001000010;
#10000;
	data_in <= 24'b011101110101000001000010;
#10000;
	data_in <= 24'b011110000101000101000011;
#10000;
	data_in <= 24'b011110010101001001000011;
#10000;
	data_in <= 24'b011111100101011001000100;
#10000;
	data_in <= 24'b100000010101100101000110;
#10000;
	data_in <= 24'b100000010101100101000110;
#10000;
	data_in <= 24'b100000100101100101000010;
#10000;
	data_in <= 24'b011101100100111101000110;
#10000;
	data_in <= 24'b011101100101000001000100;
#10000;
	data_in <= 24'b011110000101000001000100;
#10000;
	data_in <= 24'b011110100101001101000101;
#10000;
	data_in <= 24'b011111010101011001000111;
#10000;
	data_in <= 24'b100000100101101001001000;
#10000;
	data_in <= 24'b100000100101101001000111;
#10000;
	data_in <= 24'b011111110101100101000001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100000100101100001000001;
#10000;
	data_in <= 24'b100000110101101100111111;
#10000;
	data_in <= 24'b100001100101110000111111;
#10000;
	data_in <= 24'b100001110101110000111011;
#10000;
	data_in <= 24'b100010000101101100111001;
#10000;
	data_in <= 24'b100001110101101000110101;
#10000;
	data_in <= 24'b100001110101100000110010;
#10000;
	data_in <= 24'b100001000101011000101101;
#10000;
	data_in <= 24'b100001100101110001000101;
#10000;
	data_in <= 24'b100001110101111101000011;
#10000;
	data_in <= 24'b100010110101111101000010;
#10000;
	data_in <= 24'b100010100101110100111100;
#10000;
	data_in <= 24'b100010000101101000111000;
#10000;
	data_in <= 24'b100010010101101000110100;
#10000;
	data_in <= 24'b100010000101011100110001;
#10000;
	data_in <= 24'b100001100101010100101101;
#10000;
	data_in <= 24'b100010000101111001000111;
#10000;
	data_in <= 24'b100010100110001001000110;
#10000;
	data_in <= 24'b100011010110000101000100;
#10000;
	data_in <= 24'b100011010110000000111111;
#10000;
	data_in <= 24'b100010110101110100111011;
#10000;
	data_in <= 24'b100011010101111000111000;
#10000;
	data_in <= 24'b100011100101110100110111;
#10000;
	data_in <= 24'b100011010101110000110100;
#10000;
	data_in <= 24'b100010000101111001000111;
#10000;
	data_in <= 24'b100010100110001001000110;
#10000;
	data_in <= 24'b100011000110001001000101;
#10000;
	data_in <= 24'b100011000110000101000000;
#10000;
	data_in <= 24'b100011000101111100111101;
#10000;
	data_in <= 24'b100011010110000000111011;
#10000;
	data_in <= 24'b100011110110000000111010;
#10000;
	data_in <= 24'b100011110110000100111000;
#10000;
	data_in <= 24'b100001110101110101000110;
#10000;
	data_in <= 24'b100010010110000101000101;
#10000;
	data_in <= 24'b100010110110000101000100;
#10000;
	data_in <= 24'b100010110110000000111111;
#10000;
	data_in <= 24'b100010110101111000111100;
#10000;
	data_in <= 24'b100010110101111000111001;
#10000;
	data_in <= 24'b100010010101110000110110;
#10000;
	data_in <= 24'b100010000101110000110011;
#10000;
	data_in <= 24'b100001000101101101000010;
#10000;
	data_in <= 24'b100001100101111001000010;
#10000;
	data_in <= 24'b100010000101111001000001;
#10000;
	data_in <= 24'b100001110101111000111101;
#10000;
	data_in <= 24'b100010010101111100111100;
#10000;
	data_in <= 24'b100010110101111100111010;
#10000;
	data_in <= 24'b100010100101110100110111;
#10000;
	data_in <= 24'b100010000101110000110011;
#10000;
	data_in <= 24'b100000110101101001000001;
#10000;
	data_in <= 24'b100000110101101100111111;
#10000;
	data_in <= 24'b100001010101101100111110;
#10000;
	data_in <= 24'b100001100101110100111100;
#10000;
	data_in <= 24'b100010010101111100111100;
#10000;
	data_in <= 24'b100010110110000100111100;
#10000;
	data_in <= 24'b100011000110000100111010;
#10000;
	data_in <= 24'b100010100110000000110110;
#10000;
	data_in <= 24'b100001010101110001000011;
#10000;
	data_in <= 24'b100001000101110000111111;
#10000;
	data_in <= 24'b100001000101101100111011;
#10000;
	data_in <= 24'b100000110101101000111001;
#10000;
	data_in <= 24'b100001110101110100111010;
#10000;
	data_in <= 24'b100010010101111100111010;
#10000;
	data_in <= 24'b100010100101111000111001;
#10000;
	data_in <= 24'b100001110101110000110101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100010000101110000110011;
#10000;
	data_in <= 24'b100001010101101100110001;
#10000;
	data_in <= 24'b100000110101100100101111;
#10000;
	data_in <= 24'b100000100101100000101110;
#10000;
	data_in <= 24'b100000010101011000101111;
#10000;
	data_in <= 24'b100000100101011100110000;
#10000;
	data_in <= 24'b100000110101100000110001;
#10000;
	data_in <= 24'b100000110101101100110001;
#10000;
	data_in <= 24'b100010000101101100110000;
#10000;
	data_in <= 24'b100001010101101000101111;
#10000;
	data_in <= 24'b100000110101100100101110;
#10000;
	data_in <= 24'b100000110101100100101110;
#10000;
	data_in <= 24'b100000110101100100101111;
#10000;
	data_in <= 24'b100000110101100000110001;
#10000;
	data_in <= 24'b100000100101100100110010;
#10000;
	data_in <= 24'b100000110101101000110011;
#10000;
	data_in <= 24'b100010100101110100110010;
#10000;
	data_in <= 24'b100010000101111000110001;
#10000;
	data_in <= 24'b100010000101110100110010;
#10000;
	data_in <= 24'b100001110101110000110001;
#10000;
	data_in <= 24'b100001100101110000110010;
#10000;
	data_in <= 24'b100001100101110000110010;
#10000;
	data_in <= 24'b100001100101101100110100;
#10000;
	data_in <= 24'b100001100101101100110100;
#10000;
	data_in <= 24'b100011000110000100110110;
#10000;
	data_in <= 24'b100011000110001000110101;
#10000;
	data_in <= 24'b100010110110000000110101;
#10000;
	data_in <= 24'b100010010101111000110011;
#10000;
	data_in <= 24'b100001110101110100110011;
#10000;
	data_in <= 24'b100001110101110100110011;
#10000;
	data_in <= 24'b100001100101101100110100;
#10000;
	data_in <= 24'b100001010101101000110011;
#10000;
	data_in <= 24'b100010110110000000110101;
#10000;
	data_in <= 24'b100011000110000100110110;
#10000;
	data_in <= 24'b100010100101111100110100;
#10000;
	data_in <= 24'b100001110101110000110001;
#10000;
	data_in <= 24'b100001010101101100110001;
#10000;
	data_in <= 24'b100001010101101100110001;
#10000;
	data_in <= 24'b100001010101101100110001;
#10000;
	data_in <= 24'b100001000101101000110000;
#10000;
	data_in <= 24'b100010100101111000110101;
#10000;
	data_in <= 24'b100010110110000000110101;
#10000;
	data_in <= 24'b100010010101111000110011;
#10000;
	data_in <= 24'b100001100101101100110000;
#10000;
	data_in <= 24'b100001010101101100110001;
#10000;
	data_in <= 24'b100001100101110000110010;
#10000;
	data_in <= 24'b100001110101110100110011;
#10000;
	data_in <= 24'b100001010101101100110001;
#10000;
	data_in <= 24'b100010010101110100110100;
#10000;
	data_in <= 24'b100010110110000000110101;
#10000;
	data_in <= 24'b100010100101111100110100;
#10000;
	data_in <= 24'b100010000101110100110010;
#10000;
	data_in <= 24'b100001100101110000110001;
#10000;
	data_in <= 24'b100010000101111000110011;
#10000;
	data_in <= 24'b100001110101110100110011;
#10000;
	data_in <= 24'b100001010101101100110001;
#10000;
	data_in <= 24'b100010000101110000110011;
#10000;
	data_in <= 24'b100010100101111100110100;
#10000;
	data_in <= 24'b100010100101111100110100;
#10000;
	data_in <= 24'b100010000101110100110010;
#10000;
	data_in <= 24'b100001010101101100110000;
#10000;
	data_in <= 24'b100001100101110000110001;
#10000;
	data_in <= 24'b100001000101101000110000;
#10000;
	data_in <= 24'b100000010101011100101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011111110101010100101011;
#10000;
	data_in <= 24'b011111010101001100101001;
#10000;
	data_in <= 24'b011111000101001000101000;
#10000;
	data_in <= 24'b011111010101001100101000;
#10000;
	data_in <= 24'b011111010101001000100111;
#10000;
	data_in <= 24'b011110100101000000100011;
#10000;
	data_in <= 24'b011110010100111100100010;
#10000;
	data_in <= 24'b011110100101000000100011;
#10000;
	data_in <= 24'b011111100101010100101110;
#10000;
	data_in <= 24'b011110100101000100101010;
#10000;
	data_in <= 24'b011110010100111100100101;
#10000;
	data_in <= 24'b011110010100111100100100;
#10000;
	data_in <= 24'b011110110101000000100101;
#10000;
	data_in <= 24'b011110100101000000100011;
#10000;
	data_in <= 24'b011110000100111000011111;
#10000;
	data_in <= 24'b011101110100110100011110;
#10000;
	data_in <= 24'b100001100101101100110100;
#10000;
	data_in <= 24'b100000010101011000101111;
#10000;
	data_in <= 24'b011111000101001000101000;
#10000;
	data_in <= 24'b011110110101000100100110;
#10000;
	data_in <= 24'b011111100101001100101000;
#10000;
	data_in <= 24'b011111100101010000100111;
#10000;
	data_in <= 24'b011110110101000100100010;
#10000;
	data_in <= 24'b011110010100111100100000;
#10000;
	data_in <= 24'b100010010101111000110111;
#10000;
	data_in <= 24'b100001000101101000110000;
#10000;
	data_in <= 24'b100000000101011000101100;
#10000;
	data_in <= 24'b011111110101010100101010;
#10000;
	data_in <= 24'b100000000101010100101010;
#10000;
	data_in <= 24'b100000000101011000101001;
#10000;
	data_in <= 24'b011111010101001100100110;
#10000;
	data_in <= 24'b011110110101000100100010;
#10000;
	data_in <= 24'b100001000101101000110000;
#10000;
	data_in <= 24'b100000110101100100101111;
#10000;
	data_in <= 24'b100000010101011100101101;
#10000;
	data_in <= 24'b011111100101010000101001;
#10000;
	data_in <= 24'b011111010101001000100111;
#10000;
	data_in <= 24'b011111000101001000100101;
#10000;
	data_in <= 24'b011110100101000000100011;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b100000100101100000101110;
#10000;
	data_in <= 24'b100000110101100100101111;
#10000;
	data_in <= 24'b100000100101100000101101;
#10000;
	data_in <= 24'b011111110101010100101010;
#10000;
	data_in <= 24'b011111000101000100100110;
#10000;
	data_in <= 24'b011110100100111100100100;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b100000110101100100101111;
#10000;
	data_in <= 24'b100001000101101000110000;
#10000;
	data_in <= 24'b100000110101100100101111;
#10000;
	data_in <= 24'b011111110101010100101011;
#10000;
	data_in <= 24'b011110100101000000100101;
#10000;
	data_in <= 24'b011110010100111100100100;
#10000;
	data_in <= 24'b011110010100111100100100;
#10000;
	data_in <= 24'b011110000100111000100011;
#10000;
	data_in <= 24'b100000100101100000101110;
#10000;
	data_in <= 24'b100000110101100100101111;
#10000;
	data_in <= 24'b100000000101011000101100;
#10000;
	data_in <= 24'b011110110101000100100111;
#10000;
	data_in <= 24'b011110000100111000100100;
#10000;
	data_in <= 24'b011101110100110100100010;
#10000;
	data_in <= 24'b011101110100110100100011;
#10000;
	data_in <= 24'b011101100100110000100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011111000101001000100101;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011101010100101100011110;
#10000;
	data_in <= 24'b011101010100101100011110;
#10000;
	data_in <= 24'b011101100100110000011111;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011101010100101100011110;
#10000;
	data_in <= 24'b011100110100100100011100;
#10000;
	data_in <= 24'b011110010100111100100010;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011101010100101100011110;
#10000;
	data_in <= 24'b011101100100110000011111;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011110000100110100100010;
#10000;
	data_in <= 24'b011101100100101100100000;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011110010100111100100010;
#10000;
	data_in <= 24'b011110010100111100100010;
#10000;
	data_in <= 24'b011110010100111100100010;
#10000;
	data_in <= 24'b011110010100111100100010;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011110010100111100100010;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011110000100111000100001;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011101100100110000011111;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011101110100110100100000;
#10000;
	data_in <= 24'b011101100100110000011111;
#10000;
	data_in <= 24'b011101010100101100011110;
#10000;
	data_in <= 24'b011101000100101000011101;
#10000;
	data_in <= 24'b011101000100100100011110;
#10000;
	data_in <= 24'b011101000100100100011110;
#10000;
	data_in <= 24'b011101100100110000011111;
#10000;
	data_in <= 24'b011101100100110000011111;
#10000;
	data_in <= 24'b011101100100110000011111;
#10000;
	data_in <= 24'b011101100100110000011111;
#10000;
	data_in <= 24'b011101010100101100011110;
#10000;
	data_in <= 24'b011101000100101000011101;
#10000;
	data_in <= 24'b011101000100100100011110;
#10000;
	data_in <= 24'b011101000100100100011110;
#10000;
	data_in <= 24'b011101110100111000100001;
#10000;
	data_in <= 24'b011101100100110100100000;
#10000;
	data_in <= 24'b011101010100101100100000;
#10000;
	data_in <= 24'b011101000100101000011111;
#10000;
	data_in <= 24'b011101000100101000011111;
#10000;
	data_in <= 24'b011101000100101000011111;
#10000;
	data_in <= 24'b011101000100101000100000;
#10000;
	data_in <= 24'b011101000100101000100000;
#10000;
	data_in <= 24'b011101110100110100100010;
#10000;
	data_in <= 24'b011101010100101100100000;
#10000;
	data_in <= 24'b011100110100100100011110;
#10000;
	data_in <= 24'b011100100100100000011101;
#10000;
	data_in <= 24'b011100100100100000011101;
#10000;
	data_in <= 24'b011100100100100000011110;
#10000;
	data_in <= 24'b011100100100100000011110;
#10000;
	data_in <= 24'b011100010100011100011101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011100110100011000011010;
#10000;
	data_in <= 24'b011100100100011000010111;
#10000;
	data_in <= 24'b011100010100010000011000;
#10000;
	data_in <= 24'b011100100100011000010111;
#10000;
	data_in <= 24'b011100110100011100011000;
#10000;
	data_in <= 24'b011100100100011000010111;
#10000;
	data_in <= 24'b011100000100010100010100;
#10000;
	data_in <= 24'b011011100100001100010010;
#10000;
	data_in <= 24'b011110100100110100100001;
#10000;
	data_in <= 24'b011110000100101100011111;
#10000;
	data_in <= 24'b011101100100100100011101;
#10000;
	data_in <= 24'b011101010100100000011100;
#10000;
	data_in <= 24'b011101000100100000011001;
#10000;
	data_in <= 24'b011100110100011100011000;
#10000;
	data_in <= 24'b011100010100011000010101;
#10000;
	data_in <= 24'b011011110100010000010011;
#10000;
	data_in <= 24'b011111010101000000100100;
#10000;
	data_in <= 24'b011110110100111000100010;
#10000;
	data_in <= 24'b011110010100110000100000;
#10000;
	data_in <= 24'b011110000100101100011111;
#10000;
	data_in <= 24'b011101110100101100011100;
#10000;
	data_in <= 24'b011101110100101100011100;
#10000;
	data_in <= 24'b011101010100101000011001;
#10000;
	data_in <= 24'b011101000100100100011000;
#10000;
	data_in <= 24'b011110100100110100100001;
#10000;
	data_in <= 24'b011110010100110000100000;
#10000;
	data_in <= 24'b011110000100101100011111;
#10000;
	data_in <= 24'b011101110100101000011110;
#10000;
	data_in <= 24'b011101110100101100011100;
#10000;
	data_in <= 24'b011101110100101100011100;
#10000;
	data_in <= 24'b011101100100101100011010;
#10000;
	data_in <= 24'b011101000100100100011000;
#10000;
	data_in <= 24'b011101010100101000011111;
#10000;
	data_in <= 24'b011101010100101000011111;
#10000;
	data_in <= 24'b011101000100101000011101;
#10000;
	data_in <= 24'b011100110100100100011100;
#10000;
	data_in <= 24'b011100110100100100011010;
#10000;
	data_in <= 24'b011100110100100100011010;
#10000;
	data_in <= 24'b011100000100011000010111;
#10000;
	data_in <= 24'b011011010100001100010100;
#10000;
	data_in <= 24'b011100100100011100011100;
#10000;
	data_in <= 24'b011101000100100100011110;
#10000;
	data_in <= 24'b011101000100100100011110;
#10000;
	data_in <= 24'b011100110100100100011100;
#10000;
	data_in <= 24'b011101000100101000011101;
#10000;
	data_in <= 24'b011101010100101100011100;
#10000;
	data_in <= 24'b011100110100100100011010;
#10000;
	data_in <= 24'b011011110100010100010110;
#10000;
	data_in <= 24'b011100010100011100011101;
#10000;
	data_in <= 24'b011100110100100100011110;
#10000;
	data_in <= 24'b011100110100100100011110;
#10000;
	data_in <= 24'b011100100100100100011100;
#10000;
	data_in <= 24'b011101000100101100011110;
#10000;
	data_in <= 24'b011101110100111000100001;
#10000;
	data_in <= 24'b011101100100110100100000;
#10000;
	data_in <= 24'b011100110100101000011101;
#10000;
	data_in <= 24'b011100100100100000011110;
#10000;
	data_in <= 24'b011100110100100100011111;
#10000;
	data_in <= 24'b011100100100100000011110;
#10000;
	data_in <= 24'b011011100100011100011011;
#10000;
	data_in <= 24'b011100010100011100011100;
#10000;
	data_in <= 24'b011100100100101100011111;
#10000;
	data_in <= 24'b011100110100100100011110;
#10000;
	data_in <= 24'b011011100100011100011010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001011010001101000010101;
#10000;
	data_in <= 24'b001011100001101100010110;
#10000;
	data_in <= 24'b001011110001110000010111;
#10000;
	data_in <= 24'b001100100001111100011010;
#10000;
	data_in <= 24'b001101000010000100011100;
#10000;
	data_in <= 24'b001101010010001000011101;
#10000;
	data_in <= 24'b001101100010001100011110;
#10000;
	data_in <= 24'b001101100010001100011110;
#10000;
	data_in <= 24'b001011000001100100010100;
#10000;
	data_in <= 24'b001011010001101000010101;
#10000;
	data_in <= 24'b001011110001110000010111;
#10000;
	data_in <= 24'b001100010001111000011001;
#10000;
	data_in <= 24'b001100110010000000011011;
#10000;
	data_in <= 24'b001101010010001000011101;
#10000;
	data_in <= 24'b001101100010001100011110;
#10000;
	data_in <= 24'b001101110010010000011111;
#10000;
	data_in <= 24'b001010000001100000010010;
#10000;
	data_in <= 24'b001010100001101000010100;
#10000;
	data_in <= 24'b001011000001110000010110;
#10000;
	data_in <= 24'b001011100001111000011000;
#10000;
	data_in <= 24'b001100010010000100011011;
#10000;
	data_in <= 24'b001100110010001100011101;
#10000;
	data_in <= 24'b001101000010010000011110;
#10000;
	data_in <= 24'b001101010010010100011111;
#10000;
	data_in <= 24'b001010000001100000010010;
#10000;
	data_in <= 24'b001010010001100100010011;
#10000;
	data_in <= 24'b001010110001101100010101;
#10000;
	data_in <= 24'b001011010001110100010111;
#10000;
	data_in <= 24'b001011110001111100011001;
#10000;
	data_in <= 24'b001100010010000100011011;
#10000;
	data_in <= 24'b001100110010001100011101;
#10000;
	data_in <= 24'b001101010010010100011111;
#10000;
	data_in <= 24'b001001010001011100010001;
#10000;
	data_in <= 24'b001001110001100100010011;
#10000;
	data_in <= 24'b001010010001101100010101;
#10000;
	data_in <= 24'b001010100001110000010110;
#10000;
	data_in <= 24'b001011000001111000011000;
#10000;
	data_in <= 24'b001011100010000000011010;
#10000;
	data_in <= 24'b001100000010001000011100;
#10000;
	data_in <= 24'b001100100010010000011110;
#10000;
	data_in <= 24'b001001000001011000010000;
#10000;
	data_in <= 24'b001001100001100000010010;
#10000;
	data_in <= 24'b001010000001101000010100;
#10000;
	data_in <= 24'b001010100001110000010110;
#10000;
	data_in <= 24'b001010110001110100010111;
#10000;
	data_in <= 24'b001011000001111000011000;
#10000;
	data_in <= 24'b001011110010000100011011;
#10000;
	data_in <= 24'b001100010010001100011101;
#10000;
	data_in <= 24'b001000010001010100001111;
#10000;
	data_in <= 24'b001000110001011100010001;
#10000;
	data_in <= 24'b001001010001100100010011;
#10000;
	data_in <= 24'b001001110001101100010101;
#10000;
	data_in <= 24'b001010000001110000010110;
#10000;
	data_in <= 24'b001010100001111000011000;
#10000;
	data_in <= 24'b001011010010000100011101;
#10000;
	data_in <= 24'b001011110010001100011111;
#10000;
	data_in <= 24'b000111010001010000010001;
#10000;
	data_in <= 24'b001000010001011000010010;
#10000;
	data_in <= 24'b001001000001100100010001;
#10000;
	data_in <= 24'b001001100001101100010011;
#10000;
	data_in <= 24'b001010100001101100011000;
#10000;
	data_in <= 24'b001010100001111000011010;
#10000;
	data_in <= 24'b001011010010000100011101;
#10000;
	data_in <= 24'b001100100010010000011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001110000010011000011111;
#10000;
	data_in <= 24'b001110110010100000100001;
#10000;
	data_in <= 24'b001111010010101000100011;
#10000;
	data_in <= 24'b001111110010110000100101;
#10000;
	data_in <= 24'b010000000010110100100110;
#10000;
	data_in <= 24'b010000000010110100100110;
#10000;
	data_in <= 24'b010000000010110100100110;
#10000;
	data_in <= 24'b010000110010111000100110;
#10000;
	data_in <= 24'b001110010010011100100000;
#10000;
	data_in <= 24'b001110100010100000100001;
#10000;
	data_in <= 24'b001111000010101000100011;
#10000;
	data_in <= 24'b001111010010101100100100;
#10000;
	data_in <= 24'b010000000010110100100110;
#10000;
	data_in <= 24'b010000000010111000100111;
#10000;
	data_in <= 24'b010000100010111100101000;
#10000;
	data_in <= 24'b010000110011000000101001;
#10000;
	data_in <= 24'b001101110010011100100001;
#10000;
	data_in <= 24'b001110000010100000100010;
#10000;
	data_in <= 24'b001110010010100100100011;
#10000;
	data_in <= 24'b001110110010101100100101;
#10000;
	data_in <= 24'b001111100010101100100110;
#10000;
	data_in <= 24'b001111110010111100101001;
#10000;
	data_in <= 24'b010000110011000000101011;
#10000;
	data_in <= 24'b010001010011001100101100;
#10000;
	data_in <= 24'b001101100010011000100000;
#10000;
	data_in <= 24'b001110000010100000100010;
#10000;
	data_in <= 24'b001110010010100100100011;
#10000;
	data_in <= 24'b001110110010101100100101;
#10000;
	data_in <= 24'b001111010010110100100111;
#10000;
	data_in <= 24'b001111110010111100101001;
#10000;
	data_in <= 24'b010000100011001000101100;
#10000;
	data_in <= 24'b010001000011010000101110;
#10000;
	data_in <= 24'b001100110010010100011111;
#10000;
	data_in <= 24'b001101010010011100100001;
#10000;
	data_in <= 24'b001101110010100000100101;
#10000;
	data_in <= 24'b001110010010101000100111;
#10000;
	data_in <= 24'b001111000010110100101010;
#10000;
	data_in <= 24'b001111100010111100101100;
#10000;
	data_in <= 24'b010000000011000100101110;
#10000;
	data_in <= 24'b010000100011001100110000;
#10000;
	data_in <= 24'b001100110010010100011111;
#10000;
	data_in <= 24'b001101010010011100100001;
#10000;
	data_in <= 24'b001101110010100000100101;
#10000;
	data_in <= 24'b001110100010101100101000;
#10000;
	data_in <= 24'b001111010010111000101011;
#10000;
	data_in <= 24'b001111010011000100101101;
#10000;
	data_in <= 24'b010000000011010000110000;
#10000;
	data_in <= 24'b010000100011011000110010;
#10000;
	data_in <= 24'b001100100010011000100010;
#10000;
	data_in <= 24'b001100110010011100100011;
#10000;
	data_in <= 24'b001101100010101000100110;
#10000;
	data_in <= 24'b001110000010110000101000;
#10000;
	data_in <= 24'b001111000011000000101100;
#10000;
	data_in <= 24'b010000000011010000110000;
#10000;
	data_in <= 24'b010001000011100000110100;
#10000;
	data_in <= 24'b010001010011101000110110;
#10000;
	data_in <= 24'b001101010010100000100000;
#10000;
	data_in <= 24'b001101100010101000100000;
#10000;
	data_in <= 24'b001110000010110000100010;
#10000;
	data_in <= 24'b001110000010110100100101;
#10000;
	data_in <= 24'b001110110011000000101100;
#10000;
	data_in <= 24'b001111110011011000110011;
#10000;
	data_in <= 24'b010001000011101100110111;
#10000;
	data_in <= 24'b010001110011111000111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010001000011000000100101;
#10000;
	data_in <= 24'b010001000011000000100101;
#10000;
	data_in <= 24'b010001110011001000101010;
#10000;
	data_in <= 24'b010011000011011100101111;
#10000;
	data_in <= 24'b010011100011100000110010;
#10000;
	data_in <= 24'b010011100011100000110010;
#10000;
	data_in <= 24'b010011100011100000110010;
#10000;
	data_in <= 24'b010100000011101000110100;
#10000;
	data_in <= 24'b010001110011010000101100;
#10000;
	data_in <= 24'b010001100011001100101011;
#10000;
	data_in <= 24'b010010000011001100101011;
#10000;
	data_in <= 24'b010001110011010000101101;
#10000;
	data_in <= 24'b010010100011010000101110;
#10000;
	data_in <= 24'b010010000011010100101110;
#10000;
	data_in <= 24'b010010110011010100101111;
#10000;
	data_in <= 24'b010011010011011100110010;
#10000;
	data_in <= 24'b010001010011001100101100;
#10000;
	data_in <= 24'b010001010011001100101100;
#10000;
	data_in <= 24'b010001110011010000101101;
#10000;
	data_in <= 24'b010001110011010000101111;
#10000;
	data_in <= 24'b010010000011010000101111;
#10000;
	data_in <= 24'b010001110011010000101111;
#10000;
	data_in <= 24'b010010100011011000110001;
#10000;
	data_in <= 24'b010011000011011100110101;
#10000;
	data_in <= 24'b010000100011001000101100;
#10000;
	data_in <= 24'b010001000011010000101110;
#10000;
	data_in <= 24'b010001110011011100110001;
#10000;
	data_in <= 24'b010010010011100100110011;
#10000;
	data_in <= 24'b010010010011100100110011;
#10000;
	data_in <= 24'b010010000011011100110100;
#10000;
	data_in <= 24'b010010010011100000110101;
#10000;
	data_in <= 24'b010010010011100000110101;
#10000;
	data_in <= 24'b010001000011010100110010;
#10000;
	data_in <= 24'b010001100011011100110100;
#10000;
	data_in <= 24'b010010010011101000110111;
#10000;
	data_in <= 24'b010010100011101100111000;
#10000;
	data_in <= 24'b010010100011101100111000;
#10000;
	data_in <= 24'b010010010011101000111000;
#10000;
	data_in <= 24'b010010000011100100110111;
#10000;
	data_in <= 24'b010001110011100000110110;
#10000;
	data_in <= 24'b010001010011101000110110;
#10000;
	data_in <= 24'b010001110011110000111000;
#10000;
	data_in <= 24'b010010010011111000111010;
#10000;
	data_in <= 24'b010010010011111000111010;
#10000;
	data_in <= 24'b010010100011111000111100;
#10000;
	data_in <= 24'b010010110011111100111101;
#10000;
	data_in <= 24'b010010100011111000111100;
#10000;
	data_in <= 24'b010010100011110100111011;
#10000;
	data_in <= 24'b010001110011111000111011;
#10000;
	data_in <= 24'b010010010100000000111101;
#10000;
	data_in <= 24'b010010110100001000111111;
#10000;
	data_in <= 24'b010011010100010001000001;
#10000;
	data_in <= 24'b010011110100011001000011;
#10000;
	data_in <= 24'b010100000100011101000100;
#10000;
	data_in <= 24'b010011100100010101000010;
#10000;
	data_in <= 24'b010011010100000100111111;
#10000;
	data_in <= 24'b010010000100001101000000;
#10000;
	data_in <= 24'b010010010100010101000100;
#10000;
	data_in <= 24'b010011010100011101001000;
#10000;
	data_in <= 24'b010011110100100101001010;
#10000;
	data_in <= 24'b010100110100101101001011;
#10000;
	data_in <= 24'b010100100100101101001000;
#10000;
	data_in <= 24'b010011010100011001000011;
#10000;
	data_in <= 24'b010001110100000000111101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010100010011100000110100;
#10000;
	data_in <= 24'b010100010011100000110100;
#10000;
	data_in <= 24'b010100100011011100110011;
#10000;
	data_in <= 24'b010100010011011000110010;
#10000;
	data_in <= 24'b010100110011011000110010;
#10000;
	data_in <= 24'b010100110011011000110001;
#10000;
	data_in <= 24'b010101000011011000110001;
#10000;
	data_in <= 24'b010101010011100000110001;
#10000;
	data_in <= 24'b010011110011100100110100;
#10000;
	data_in <= 24'b010100010011100000110100;
#10000;
	data_in <= 24'b010100000011011100110011;
#10000;
	data_in <= 24'b010100010011011000110010;
#10000;
	data_in <= 24'b010100000011010100110001;
#10000;
	data_in <= 24'b010100100011010100110001;
#10000;
	data_in <= 24'b010100100011010100110000;
#10000;
	data_in <= 24'b010100100011010100110000;
#10000;
	data_in <= 24'b010011000011011100110101;
#10000;
	data_in <= 24'b010011100011011100110101;
#10000;
	data_in <= 24'b010011010011011000110100;
#10000;
	data_in <= 24'b010011110011011000110100;
#10000;
	data_in <= 24'b010011100011010100110001;
#10000;
	data_in <= 24'b010100000011010100110001;
#10000;
	data_in <= 24'b010011110011010000110000;
#10000;
	data_in <= 24'b010011110011010100101111;
#10000;
	data_in <= 24'b010010010011011000110011;
#10000;
	data_in <= 24'b010010010011011000110011;
#10000;
	data_in <= 24'b010010100011010100110011;
#10000;
	data_in <= 24'b010010100011010100110011;
#10000;
	data_in <= 24'b010011000011011000110001;
#10000;
	data_in <= 24'b010011000011011000110001;
#10000;
	data_in <= 24'b010011100011010100110001;
#10000;
	data_in <= 24'b010011100011010100110001;
#10000;
	data_in <= 24'b010010000011011000110101;
#10000;
	data_in <= 24'b010010000011011000110101;
#10000;
	data_in <= 24'b010010010011011000110011;
#10000;
	data_in <= 24'b010010010011011000110011;
#10000;
	data_in <= 24'b010010010011010100110000;
#10000;
	data_in <= 24'b010010010011010100110000;
#10000;
	data_in <= 24'b010010110011010100110000;
#10000;
	data_in <= 24'b010010110011010100110000;
#10000;
	data_in <= 24'b010010000011101100111001;
#10000;
	data_in <= 24'b010010100011101100111001;
#10000;
	data_in <= 24'b010010000011100100110110;
#10000;
	data_in <= 24'b010010000011011100110100;
#10000;
	data_in <= 24'b010001110011011100110001;
#10000;
	data_in <= 24'b010001110011010000101111;
#10000;
	data_in <= 24'b010001110011010000101111;
#10000;
	data_in <= 24'b010010000011010000101111;
#10000;
	data_in <= 24'b010011000100000000111110;
#10000;
	data_in <= 24'b010010110011111000111100;
#10000;
	data_in <= 24'b010010010011110100111001;
#10000;
	data_in <= 24'b010010000011100100110110;
#10000;
	data_in <= 24'b010001010011011100110001;
#10000;
	data_in <= 24'b010001100011011000110000;
#10000;
	data_in <= 24'b010001100011011000110000;
#10000;
	data_in <= 24'b010001110011010000101111;
#10000;
	data_in <= 24'b010010100100001001000010;
#10000;
	data_in <= 24'b010010000100000001000000;
#10000;
	data_in <= 24'b010001110011110100111101;
#10000;
	data_in <= 24'b010001000011101100111000;
#10000;
	data_in <= 24'b010000110011011100110111;
#10000;
	data_in <= 24'b010000110011011000110100;
#10000;
	data_in <= 24'b010001010011011100110001;
#10000;
	data_in <= 24'b010010000011100000110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b010101000011100000110001;
#10000;
	data_in <= 24'b010101100011101000110011;
#10000;
	data_in <= 24'b010101110011101100110100;
#10000;
	data_in <= 24'b010110000011101100110100;
#10000;
	data_in <= 24'b010110100011101000110100;
#10000;
	data_in <= 24'b010110110011101100110101;
#10000;
	data_in <= 24'b011000000011111000111000;
#10000;
	data_in <= 24'b011000100100000000111010;
#10000;
	data_in <= 24'b010100000011011000110000;
#10000;
	data_in <= 24'b010100100011100000110001;
#10000;
	data_in <= 24'b010101010011100100110010;
#10000;
	data_in <= 24'b010101100011101000110011;
#10000;
	data_in <= 24'b010110000011101100110100;
#10000;
	data_in <= 24'b010110110011101100110101;
#10000;
	data_in <= 24'b011000000011111000111000;
#10000;
	data_in <= 24'b011000100100000000111010;
#10000;
	data_in <= 24'b010100010011011100110001;
#10000;
	data_in <= 24'b010011110011011100110001;
#10000;
	data_in <= 24'b010100110011100100110011;
#10000;
	data_in <= 24'b010101100011100100110100;
#10000;
	data_in <= 24'b010110000011101000110101;
#10000;
	data_in <= 24'b010110100011110000110111;
#10000;
	data_in <= 24'b010111010011110100111000;
#10000;
	data_in <= 24'b010111100011111000111001;
#10000;
	data_in <= 24'b010100000011100000110010;
#10000;
	data_in <= 24'b010100010011100100110011;
#10000;
	data_in <= 24'b010100110011100100110011;
#10000;
	data_in <= 24'b010101000011101000110100;
#10000;
	data_in <= 24'b010101110011101000110101;
#10000;
	data_in <= 24'b010110010011101100110110;
#10000;
	data_in <= 24'b010111000011110000110111;
#10000;
	data_in <= 24'b010111000011110000110111;
#10000;
	data_in <= 24'b010011110011011000110010;
#10000;
	data_in <= 24'b010100000011011100110011;
#10000;
	data_in <= 24'b010100110011100100110011;
#10000;
	data_in <= 24'b010101000011101000110100;
#10000;
	data_in <= 24'b010101110011101000110101;
#10000;
	data_in <= 24'b010101110011101000110101;
#10000;
	data_in <= 24'b010110100011101100111000;
#10000;
	data_in <= 24'b010110100011101100111000;
#10000;
	data_in <= 24'b010010100011010000101111;
#10000;
	data_in <= 24'b010011100011010100110001;
#10000;
	data_in <= 24'b010100100011100000110010;
#10000;
	data_in <= 24'b010100110011100100110011;
#10000;
	data_in <= 24'b010101010011100000110011;
#10000;
	data_in <= 24'b010101110011101000110101;
#10000;
	data_in <= 24'b010110110011110000111001;
#10000;
	data_in <= 24'b010111010011111000111011;
#10000;
	data_in <= 24'b010010100011010000101111;
#10000;
	data_in <= 24'b010011000011011000110001;
#10000;
	data_in <= 24'b010100000011011100110011;
#10000;
	data_in <= 24'b010100110011100000110100;
#10000;
	data_in <= 24'b010101010011100000110100;
#10000;
	data_in <= 24'b010101110011101000110110;
#10000;
	data_in <= 24'b010111000011111100111011;
#10000;
	data_in <= 24'b010111110100001000111110;
#10000;
	data_in <= 24'b010010010011011100110000;
#10000;
	data_in <= 24'b010011000011100100110010;
#10000;
	data_in <= 24'b010011110011101100110110;
#10000;
	data_in <= 24'b010011100011101000110101;
#10000;
	data_in <= 24'b010101000011101000110100;
#10000;
	data_in <= 24'b010101110011101100110100;
#10000;
	data_in <= 24'b010111110011111100111001;
#10000;
	data_in <= 24'b011001000100001101000000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011001100100001000111100;
#10000;
	data_in <= 24'b011001110100001100111011;
#10000;
	data_in <= 24'b011010010100010100111111;
#10000;
	data_in <= 24'b011010110100011100111111;
#10000;
	data_in <= 24'b011011110100100101000100;
#10000;
	data_in <= 24'b011011110100101101000011;
#10000;
	data_in <= 24'b011100100100110101000101;
#10000;
	data_in <= 24'b011100100100110101000101;
#10000;
	data_in <= 24'b011001010100000100111011;
#10000;
	data_in <= 24'b011001100100001000111100;
#10000;
	data_in <= 24'b011010000100010000111110;
#10000;
	data_in <= 24'b011010000100011001000000;
#10000;
	data_in <= 24'b011011000100011101000011;
#10000;
	data_in <= 24'b011011000100100101000101;
#10000;
	data_in <= 24'b011011010100101001000110;
#10000;
	data_in <= 24'b011011100100110001000110;
#10000;
	data_in <= 24'b011000110100000000111100;
#10000;
	data_in <= 24'b011001000100000100111101;
#10000;
	data_in <= 24'b011001010100001000111110;
#10000;
	data_in <= 24'b011001010100010101000000;
#10000;
	data_in <= 24'b011010010100011001000011;
#10000;
	data_in <= 24'b011010010100100001000101;
#10000;
	data_in <= 24'b011010110100101001000111;
#10000;
	data_in <= 24'b011010110100101001000111;
#10000;
	data_in <= 24'b011000010100000100111100;
#10000;
	data_in <= 24'b011000100100000100111110;
#10000;
	data_in <= 24'b011000110100001000111111;
#10000;
	data_in <= 24'b011001100100010001000100;
#10000;
	data_in <= 24'b011010000100011001000110;
#10000;
	data_in <= 24'b011010000100100101001000;
#10000;
	data_in <= 24'b011010100100101001001011;
#10000;
	data_in <= 24'b011010110100110001001011;
#10000;
	data_in <= 24'b010111100011111100111100;
#10000;
	data_in <= 24'b010111110100000000111111;
#10000;
	data_in <= 24'b011000010100001001000001;
#10000;
	data_in <= 24'b011001000100010001000101;
#10000;
	data_in <= 24'b011001100100011001000111;
#10000;
	data_in <= 24'b011010000100100101001010;
#10000;
	data_in <= 24'b011010100100101101001110;
#10000;
	data_in <= 24'b011010110100110001001111;
#10000;
	data_in <= 24'b010111100011111100111110;
#10000;
	data_in <= 24'b010111110100000000111111;
#10000;
	data_in <= 24'b011000100100001001000011;
#10000;
	data_in <= 24'b011001000100010101001000;
#10000;
	data_in <= 24'b011001110100100001001011;
#10000;
	data_in <= 24'b011001110100100101001110;
#10000;
	data_in <= 24'b011010000100101001001111;
#10000;
	data_in <= 24'b011010010100101101010000;
#10000;
	data_in <= 24'b011000010100001101000010;
#10000;
	data_in <= 24'b011000110100010001000101;
#10000;
	data_in <= 24'b011001100100011101001010;
#10000;
	data_in <= 24'b011001110100101001001101;
#10000;
	data_in <= 24'b011010010100101101010000;
#10000;
	data_in <= 24'b011010010100110101010011;
#10000;
	data_in <= 24'b011010010100110101010011;
#10000;
	data_in <= 24'b011010010100111001010010;
#10000;
	data_in <= 24'b011001110100011001001010;
#10000;
	data_in <= 24'b011010000100100001001101;
#10000;
	data_in <= 24'b011001110100101101010001;
#10000;
	data_in <= 24'b011010000100111001010100;
#10000;
	data_in <= 24'b011010100101000001010110;
#10000;
	data_in <= 24'b011010010101001001010111;
#10000;
	data_in <= 24'b011010010101000001011010;
#10000;
	data_in <= 24'b011001110101000001011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011100100100110101000101;
#10000;
	data_in <= 24'b011100110100111101000101;
#10000;
	data_in <= 24'b011101100100111101000110;
#10000;
	data_in <= 24'b011101110101000101000101;
#10000;
	data_in <= 24'b011110010101001001000011;
#10000;
	data_in <= 24'b011110100101010001000010;
#10000;
	data_in <= 24'b011111010101010101000010;
#10000;
	data_in <= 24'b011111100101100001000000;
#10000;
	data_in <= 24'b011100100100111001001000;
#10000;
	data_in <= 24'b011100110100111101000111;
#10000;
	data_in <= 24'b011101000101000001001000;
#10000;
	data_in <= 24'b011101010101001001000101;
#10000;
	data_in <= 24'b011101110101001001000100;
#10000;
	data_in <= 24'b011110010101001101000001;
#10000;
	data_in <= 24'b011111000101010001000001;
#10000;
	data_in <= 24'b011111000101011000111110;
#10000;
	data_in <= 24'b011011110100110001001000;
#10000;
	data_in <= 24'b011100010100111101001001;
#10000;
	data_in <= 24'b011100100101000101001000;
#10000;
	data_in <= 24'b011101010101001001001000;
#10000;
	data_in <= 24'b011101110101000101000101;
#10000;
	data_in <= 24'b011110010101001001000011;
#10000;
	data_in <= 24'b011110110101001101000000;
#10000;
	data_in <= 24'b011110110101010100111101;
#10000;
	data_in <= 24'b011010100100101101001000;
#10000;
	data_in <= 24'b011011010100110101001000;
#10000;
	data_in <= 24'b011011110100111101001001;
#10000;
	data_in <= 24'b011100100101001001000111;
#10000;
	data_in <= 24'b011101010101001001000101;
#10000;
	data_in <= 24'b011101110101001101000011;
#10000;
	data_in <= 24'b011110010101010001000000;
#10000;
	data_in <= 24'b011110110101010100111101;
#10000;
	data_in <= 24'b011010100100110001001011;
#10000;
	data_in <= 24'b011011000100110101001010;
#10000;
	data_in <= 24'b011100000101000001001010;
#10000;
	data_in <= 24'b011100100101000101001000;
#10000;
	data_in <= 24'b011101010101001001000101;
#10000;
	data_in <= 24'b011101110101001101000011;
#10000;
	data_in <= 24'b011110010101010001000000;
#10000;
	data_in <= 24'b011110110101010100111101;
#10000;
	data_in <= 24'b011010110100111101001111;
#10000;
	data_in <= 24'b011011100101000101001101;
#10000;
	data_in <= 24'b011011110101000101001100;
#10000;
	data_in <= 24'b011100010101001001001001;
#10000;
	data_in <= 24'b011101000101001001000101;
#10000;
	data_in <= 24'b011101000101001001000010;
#10000;
	data_in <= 24'b011110000101001100111111;
#10000;
	data_in <= 24'b011110100101010000111100;
#10000;
	data_in <= 24'b011011100101001001010010;
#10000;
	data_in <= 24'b011100000101001101001111;
#10000;
	data_in <= 24'b011100010101001101001110;
#10000;
	data_in <= 24'b011100100101001001001100;
#10000;
	data_in <= 24'b011101010101001001001000;
#10000;
	data_in <= 24'b011101010101001001000100;
#10000;
	data_in <= 24'b011110010101010001000000;
#10000;
	data_in <= 24'b011111000101011000111110;
#10000;
	data_in <= 24'b011001010101001001010101;
#10000;
	data_in <= 24'b011001110101001001010100;
#10000;
	data_in <= 24'b011011100101001001010001;
#10000;
	data_in <= 24'b011100100101000101001110;
#10000;
	data_in <= 24'b011101010101000101001001;
#10000;
	data_in <= 24'b011101110101010001000111;
#10000;
	data_in <= 24'b011110100101011001000110;
#10000;
	data_in <= 24'b011110110101100101000010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100000100101100101000000;
#10000;
	data_in <= 24'b100000010101100100111100;
#10000;
	data_in <= 24'b100000110101101000111010;
#10000;
	data_in <= 24'b100000100101100100111000;
#10000;
	data_in <= 24'b100000100101101000110111;
#10000;
	data_in <= 24'b100001000101110100110111;
#10000;
	data_in <= 24'b100010000101111000111001;
#10000;
	data_in <= 24'b100010100110000100111010;
#10000;
	data_in <= 24'b011111110101011000111101;
#10000;
	data_in <= 24'b011111110101011100111010;
#10000;
	data_in <= 24'b100000010101100000111000;
#10000;
	data_in <= 24'b100000010101100000110111;
#10000;
	data_in <= 24'b100000010101100100110110;
#10000;
	data_in <= 24'b100000100101101000110111;
#10000;
	data_in <= 24'b100001100101110000110111;
#10000;
	data_in <= 24'b100010000101111000111001;
#10000;
	data_in <= 24'b011111010101010000111011;
#10000;
	data_in <= 24'b011111100101011000111001;
#10000;
	data_in <= 24'b100000010101100000111000;
#10000;
	data_in <= 24'b100000010101100000110111;
#10000;
	data_in <= 24'b100000010101100100110110;
#10000;
	data_in <= 24'b100000100101101000110111;
#10000;
	data_in <= 24'b100001000101110100110111;
#10000;
	data_in <= 24'b100001010101111000111000;
#10000;
	data_in <= 24'b011111100101010100111100;
#10000;
	data_in <= 24'b011111110101011100111010;
#10000;
	data_in <= 24'b100000110101101000111010;
#10000;
	data_in <= 24'b100000110101101000111001;
#10000;
	data_in <= 24'b100000110101101100111000;
#10000;
	data_in <= 24'b100000110101101100111000;
#10000;
	data_in <= 24'b100001000101110100110111;
#10000;
	data_in <= 24'b100001010101111000111000;
#10000;
	data_in <= 24'b011111110101011000111101;
#10000;
	data_in <= 24'b100000000101100000111011;
#10000;
	data_in <= 24'b100001000101101100111011;
#10000;
	data_in <= 24'b100001000101101100111010;
#10000;
	data_in <= 24'b100001000101110000111001;
#10000;
	data_in <= 24'b100001000101110000111001;
#10000;
	data_in <= 24'b100001000101110100110111;
#10000;
	data_in <= 24'b100001000101110100110111;
#10000;
	data_in <= 24'b011111100101011000111101;
#10000;
	data_in <= 24'b100000000101100000111011;
#10000;
	data_in <= 24'b100001000101101100111011;
#10000;
	data_in <= 24'b100001010101110000111011;
#10000;
	data_in <= 24'b100001010101110100111010;
#10000;
	data_in <= 24'b100001010101110100111010;
#10000;
	data_in <= 24'b100001010101111000111000;
#10000;
	data_in <= 24'b100001010101111000111000;
#10000;
	data_in <= 24'b011111110101011100111110;
#10000;
	data_in <= 24'b100000100101101000111101;
#10000;
	data_in <= 24'b100001100101110100111101;
#10000;
	data_in <= 24'b100001110101111000111101;
#10000;
	data_in <= 24'b100010100110000000111101;
#10000;
	data_in <= 24'b100010110110000100111110;
#10000;
	data_in <= 24'b100010110110000100111110;
#10000;
	data_in <= 24'b100011000110001000111111;
#10000;
	data_in <= 24'b011111010101100101000001;
#10000;
	data_in <= 24'b100000010101110001000000;
#10000;
	data_in <= 24'b100000110101111101000001;
#10000;
	data_in <= 24'b100001110110000101000001;
#10000;
	data_in <= 24'b100010010110010001000010;
#10000;
	data_in <= 24'b100010110110010101000011;
#10000;
	data_in <= 24'b100011100110011001000011;
#10000;
	data_in <= 24'b100011110110011101000100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100001110101110100110011;
#10000;
	data_in <= 24'b100001100101110000110010;
#10000;
	data_in <= 24'b100001100101110000110001;
#10000;
	data_in <= 24'b100001100101110000110001;
#10000;
	data_in <= 24'b100001100101110000110001;
#10000;
	data_in <= 24'b100001000101101000101111;
#10000;
	data_in <= 24'b100000100101100000101101;
#10000;
	data_in <= 24'b100000000101011000101011;
#10000;
	data_in <= 24'b100001100101101100110100;
#10000;
	data_in <= 24'b100001010101101100110001;
#10000;
	data_in <= 24'b100001000101101000110000;
#10000;
	data_in <= 24'b100001000101101000101111;
#10000;
	data_in <= 24'b100001000101101000101111;
#10000;
	data_in <= 24'b100000110101100100101110;
#10000;
	data_in <= 24'b100000000101011000101011;
#10000;
	data_in <= 24'b011111100101010000101001;
#10000;
	data_in <= 24'b100001010101110000110101;
#10000;
	data_in <= 24'b100001000101110000110010;
#10000;
	data_in <= 24'b100000100101101000110000;
#10000;
	data_in <= 24'b100000100101101000110000;
#10000;
	data_in <= 24'b100000010101100100101111;
#10000;
	data_in <= 24'b100000000101100000101110;
#10000;
	data_in <= 24'b011111100101011000101100;
#10000;
	data_in <= 24'b011111000101010000101010;
#10000;
	data_in <= 24'b100001110101111000110111;
#10000;
	data_in <= 24'b100001010101110000110101;
#10000;
	data_in <= 24'b100001000101101100110100;
#10000;
	data_in <= 24'b100000110101101100110001;
#10000;
	data_in <= 24'b100000100101101000110000;
#10000;
	data_in <= 24'b100000010101100100101111;
#10000;
	data_in <= 24'b011111110101011100101101;
#10000;
	data_in <= 24'b011111010101010100101011;
#10000;
	data_in <= 24'b100001100101111100111001;
#10000;
	data_in <= 24'b100001000101110100110110;
#10000;
	data_in <= 24'b100000110101110000110101;
#10000;
	data_in <= 24'b100000100101101100110100;
#10000;
	data_in <= 24'b100000110101101100110001;
#10000;
	data_in <= 24'b100000100101101000110000;
#10000;
	data_in <= 24'b011111110101011100101101;
#10000;
	data_in <= 24'b011111010101010100101011;
#10000;
	data_in <= 24'b100001110110000000111010;
#10000;
	data_in <= 24'b100001100101111100111001;
#10000;
	data_in <= 24'b100001010101111000110111;
#10000;
	data_in <= 24'b100001000101110100110110;
#10000;
	data_in <= 24'b100001100101110100110110;
#10000;
	data_in <= 24'b100001000101110000110010;
#10000;
	data_in <= 24'b100000010101100100101111;
#10000;
	data_in <= 24'b011111110101011100101101;
#10000;
	data_in <= 24'b100010110110010000111110;
#10000;
	data_in <= 24'b100010100110001100111101;
#10000;
	data_in <= 24'b100010010110001000111100;
#10000;
	data_in <= 24'b100010010110001000111011;
#10000;
	data_in <= 24'b100010010110001000111011;
#10000;
	data_in <= 24'b100001110110000000111001;
#10000;
	data_in <= 24'b100001000101111000110100;
#10000;
	data_in <= 24'b100000010101101100110001;
#10000;
	data_in <= 24'b100011110110100001000010;
#10000;
	data_in <= 24'b100011110110100001000001;
#10000;
	data_in <= 24'b100011110110100001000010;
#10000;
	data_in <= 24'b100100010110100001000001;
#10000;
	data_in <= 24'b100100010110100001000001;
#10000;
	data_in <= 24'b100011100110011000111100;
#10000;
	data_in <= 24'b100010110110001100111001;
#10000;
	data_in <= 24'b100010000110000000110110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011111110101010100101011;
#10000;
	data_in <= 24'b011111110101010100101011;
#10000;
	data_in <= 24'b011111000101010000101010;
#10000;
	data_in <= 24'b011110100101001000101000;
#10000;
	data_in <= 24'b011101110100111100100101;
#10000;
	data_in <= 24'b011101010100110100100011;
#10000;
	data_in <= 24'b011100110100101000100011;
#10000;
	data_in <= 24'b011100110100101100100001;
#10000;
	data_in <= 24'b011110110101000100100111;
#10000;
	data_in <= 24'b011110100101001000101000;
#10000;
	data_in <= 24'b011110010101000100100111;
#10000;
	data_in <= 24'b011110000100111100101000;
#10000;
	data_in <= 24'b011101100100110100100110;
#10000;
	data_in <= 24'b011101000100101100100100;
#10000;
	data_in <= 24'b011100110100100100100100;
#10000;
	data_in <= 24'b011100010100101000100011;
#10000;
	data_in <= 24'b011110100101001000101000;
#10000;
	data_in <= 24'b011110100101001000101000;
#10000;
	data_in <= 24'b011110010101000000101001;
#10000;
	data_in <= 24'b011101010100111000100111;
#10000;
	data_in <= 24'b011100110100110000100110;
#10000;
	data_in <= 24'b011100000100100100100011;
#10000;
	data_in <= 24'b011011110100011100100100;
#10000;
	data_in <= 24'b011011010100100000100010;
#10000;
	data_in <= 24'b011111000101010000101010;
#10000;
	data_in <= 24'b011110010101001100101001;
#10000;
	data_in <= 24'b011101110101000000101001;
#10000;
	data_in <= 24'b011101010100111000101000;
#10000;
	data_in <= 24'b011100110100101100101000;
#10000;
	data_in <= 24'b011011110100100100100110;
#10000;
	data_in <= 24'b011011010100011100100100;
#10000;
	data_in <= 24'b011011010100011100100100;
#10000;
	data_in <= 24'b011101110101000000101001;
#10000;
	data_in <= 24'b011101110101000000101001;
#10000;
	data_in <= 24'b011101010100111000101000;
#10000;
	data_in <= 24'b011100100100110100100111;
#10000;
	data_in <= 24'b011100010100101100101000;
#10000;
	data_in <= 24'b011100000100101000101000;
#10000;
	data_in <= 24'b011100000100101000101000;
#10000;
	data_in <= 24'b011011110100101000101000;
#10000;
	data_in <= 24'b011110100101001100101100;
#10000;
	data_in <= 24'b011110000101000100101010;
#10000;
	data_in <= 24'b011101000100111100101001;
#10000;
	data_in <= 24'b011100010100101100101000;
#10000;
	data_in <= 24'b011100000100101000101000;
#10000;
	data_in <= 24'b011011100100100100100111;
#10000;
	data_in <= 24'b011011010100011100100111;
#10000;
	data_in <= 24'b011011000100011000100110;
#10000;
	data_in <= 24'b011111100101011100110000;
#10000;
	data_in <= 24'b011110110101010000101101;
#10000;
	data_in <= 24'b011101010101000000101010;
#10000;
	data_in <= 24'b011100100100110000101001;
#10000;
	data_in <= 24'b011011100100100100100111;
#10000;
	data_in <= 24'b011011000100011000100110;
#10000;
	data_in <= 24'b011010100100010000100110;
#10000;
	data_in <= 24'b011001110100001100100101;
#10000;
	data_in <= 24'b100000000101011100110000;
#10000;
	data_in <= 24'b011111100101010000101111;
#10000;
	data_in <= 24'b011110000101000000101101;
#10000;
	data_in <= 24'b011100100100110000101010;
#10000;
	data_in <= 24'b011100000100100100101001;
#10000;
	data_in <= 24'b011011010100011100101001;
#10000;
	data_in <= 24'b011010110100010100100111;
#10000;
	data_in <= 24'b011010000100010000100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011100000100100000011110;
#10000;
	data_in <= 24'b011011110100011100011101;
#10000;
	data_in <= 24'b011011110100011100011101;
#10000;
	data_in <= 24'b011100000100100000011110;
#10000;
	data_in <= 24'b011100000100100000011110;
#10000;
	data_in <= 24'b011011100100010100011110;
#10000;
	data_in <= 24'b011011100100010100011110;
#10000;
	data_in <= 24'b011011110100011000011111;
#10000;
	data_in <= 24'b011011110100011000011111;
#10000;
	data_in <= 24'b011011010100011000011111;
#10000;
	data_in <= 24'b011011110100011000011111;
#10000;
	data_in <= 24'b011011100100011100100000;
#10000;
	data_in <= 24'b011100000100011100100000;
#10000;
	data_in <= 24'b011011010100011000100000;
#10000;
	data_in <= 24'b011011110100010100100000;
#10000;
	data_in <= 24'b011011110100100000100010;
#10000;
	data_in <= 24'b011010110100010000011110;
#10000;
	data_in <= 24'b011010000100001100011101;
#10000;
	data_in <= 24'b011010110100010000011110;
#10000;
	data_in <= 24'b011010100100010100011111;
#10000;
	data_in <= 24'b011011000100010100011111;
#10000;
	data_in <= 24'b011010010100001100100000;
#10000;
	data_in <= 24'b011011000100010000100001;
#10000;
	data_in <= 24'b011011000100011000100011;
#10000;
	data_in <= 24'b011010100100010000100001;
#10000;
	data_in <= 24'b011010000100001000011111;
#10000;
	data_in <= 24'b011001110100000100011110;
#10000;
	data_in <= 24'b011010000100001000100000;
#10000;
	data_in <= 24'b011010010100001100100001;
#10000;
	data_in <= 24'b011010000100001000100000;
#10000;
	data_in <= 24'b011010000100001000100000;
#10000;
	data_in <= 24'b011010000100001100100001;
#10000;
	data_in <= 24'b011011100100100100100111;
#10000;
	data_in <= 24'b011010010100010000100010;
#10000;
	data_in <= 24'b011001100100000100011111;
#10000;
	data_in <= 24'b011001110100000100100001;
#10000;
	data_in <= 24'b011010010100001100100011;
#10000;
	data_in <= 24'b011010000100001000100010;
#10000;
	data_in <= 24'b011001110100000100100001;
#10000;
	data_in <= 24'b011000110100000000011111;
#10000;
	data_in <= 24'b011011100100100000101000;
#10000;
	data_in <= 24'b011010010100001100100011;
#10000;
	data_in <= 24'b011001010011111100011111;
#10000;
	data_in <= 24'b011001010011111100011111;
#10000;
	data_in <= 24'b011001110100000100100011;
#10000;
	data_in <= 24'b011001010100000100100011;
#10000;
	data_in <= 24'b011000110011111100100001;
#10000;
	data_in <= 24'b011000100011111000100000;
#10000;
	data_in <= 24'b011010000100010000100110;
#10000;
	data_in <= 24'b011001000100000000100010;
#10000;
	data_in <= 24'b011000100011111000100000;
#10000;
	data_in <= 24'b011000100011111000100000;
#10000;
	data_in <= 24'b011000110011111000100010;
#10000;
	data_in <= 24'b011000100011110100100001;
#10000;
	data_in <= 24'b011000100011110100100001;
#10000;
	data_in <= 24'b011000010011111100100010;
#10000;
	data_in <= 24'b011001010100000100100011;
#10000;
	data_in <= 24'b011001000100000000100010;
#10000;
	data_in <= 24'b011000110011111100100001;
#10000;
	data_in <= 24'b011000110011111100100001;
#10000;
	data_in <= 24'b011000100011110100100001;
#10000;
	data_in <= 24'b011000000011111000100001;
#10000;
	data_in <= 24'b011000100011111100100101;
#10000;
	data_in <= 24'b011000100100000100100111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011010100010000011101;
#10000;
	data_in <= 24'b011011100100010100011110;
#10000;
	data_in <= 24'b011011100100010100011110;
#10000;
	data_in <= 24'b011011000100011000011100;
#10000;
	data_in <= 24'b011011110100011100011101;
#10000;
	data_in <= 24'b011011100100100000011110;
#10000;
	data_in <= 24'b011011110100011100011101;
#10000;
	data_in <= 24'b011010110100011000011010;
#10000;
	data_in <= 24'b011011010100001100011110;
#10000;
	data_in <= 24'b011011000100010100011111;
#10000;
	data_in <= 24'b011010110100010000011110;
#10000;
	data_in <= 24'b011010110100010000011110;
#10000;
	data_in <= 24'b011011000100010100011111;
#10000;
	data_in <= 24'b011011100100011100100000;
#10000;
	data_in <= 24'b011011010100011000011111;
#10000;
	data_in <= 24'b011010100100011000011110;
#10000;
	data_in <= 24'b011011100100011000100011;
#10000;
	data_in <= 24'b011011000100011000100011;
#10000;
	data_in <= 24'b011010100100010000100001;
#10000;
	data_in <= 24'b011010000100001000011111;
#10000;
	data_in <= 24'b011010000100001000011111;
#10000;
	data_in <= 24'b011010010100010000011110;
#10000;
	data_in <= 24'b011010010100010000011110;
#10000;
	data_in <= 24'b011001110100001100011101;
#10000;
	data_in <= 24'b011010100100001100100011;
#10000;
	data_in <= 24'b011010100100010100100011;
#10000;
	data_in <= 24'b011010100100001100100011;
#10000;
	data_in <= 24'b011001110100001000100000;
#10000;
	data_in <= 24'b011001110100000100011111;
#10000;
	data_in <= 24'b011001110100001000100000;
#10000;
	data_in <= 24'b011010000100001100100001;
#10000;
	data_in <= 24'b011001110100001000100000;
#10000;
	data_in <= 24'b011001000011111000100000;
#10000;
	data_in <= 24'b011000110100000000011111;
#10000;
	data_in <= 24'b011001100100000000100010;
#10000;
	data_in <= 24'b011001000100000100100000;
#10000;
	data_in <= 24'b011001100100000000100000;
#10000;
	data_in <= 24'b011001100100001100100010;
#10000;
	data_in <= 24'b011001100100001100100010;
#10000;
	data_in <= 24'b011001100100001100100010;
#10000;
	data_in <= 24'b011000100011110100100001;
#10000;
	data_in <= 24'b011001000100000000100010;
#10000;
	data_in <= 24'b011001010100000000100100;
#10000;
	data_in <= 24'b011001000100000000100010;
#10000;
	data_in <= 24'b011001000100000000100010;
#10000;
	data_in <= 24'b011001010100000100100011;
#10000;
	data_in <= 24'b011001100100001000100100;
#10000;
	data_in <= 24'b011001010100000100100011;
#10000;
	data_in <= 24'b011001000100000100100111;
#10000;
	data_in <= 24'b011001010100001100100110;
#10000;
	data_in <= 24'b011001010100001000101000;
#10000;
	data_in <= 24'b011001000100001000100101;
#10000;
	data_in <= 24'b011001000100001000100101;
#10000;
	data_in <= 24'b011001010100001100100110;
#10000;
	data_in <= 24'b011001110100010100101000;
#10000;
	data_in <= 24'b011001110100010100101000;
#10000;
	data_in <= 24'b011000010100000000100110;
#10000;
	data_in <= 24'b011000110100000100101001;
#10000;
	data_in <= 24'b011000100100001100101010;
#10000;
	data_in <= 24'b011000100100001100101010;
#10000;
	data_in <= 24'b011000110100010000101011;
#10000;
	data_in <= 24'b011001100100100000101111;
#10000;
	data_in <= 24'b011010010100101100110010;
#10000;
	data_in <= 24'b011010110100110100110100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000111010001100000011010;
#10000;
	data_in <= 24'b000111100001100100010110;
#10000;
	data_in <= 24'b001010010001111100010101;
#10000;
	data_in <= 24'b001010010001110100010011;
#10000;
	data_in <= 24'b001011010001101100011010;
#10000;
	data_in <= 24'b001011110001111100100000;
#10000;
	data_in <= 24'b001010110001110000011001;
#10000;
	data_in <= 24'b001010100001101100010010;
#10000;
	data_in <= 24'b000011010000110000010000;
#10000;
	data_in <= 24'b000100100001000000010000;
#10000;
	data_in <= 24'b000111100001010100010001;
#10000;
	data_in <= 24'b000111100001001100001111;
#10000;
	data_in <= 24'b000111100001000000010100;
#10000;
	data_in <= 24'b001001100001100000011110;
#10000;
	data_in <= 24'b001101100010100100100111;
#10000;
	data_in <= 24'b010110110100110001000011;
#10000;
	data_in <= 24'b000001000000010100001001;
#10000;
	data_in <= 24'b000000010000000000000101;
#10000;
	data_in <= 24'b000001110000000000001001;
#10000;
	data_in <= 24'b000010110000010100010000;
#10000;
	data_in <= 24'b000001100000000100010000;
#10000;
	data_in <= 24'b000011010000011000010011;
#10000;
	data_in <= 24'b001100100010100000101110;
#10000;
	data_in <= 24'b100010110111101101110101;
#10000;
	data_in <= 24'b000001010000010100000101;
#10000;
	data_in <= 24'b000011010000110000010000;
#10000;
	data_in <= 24'b000011000000100000010100;
#10000;
	data_in <= 24'b000001110000001100010110;
#10000;
	data_in <= 24'b000010010000101100011101;
#10000;
	data_in <= 24'b000101100001011100100101;
#10000;
	data_in <= 24'b001000010001110100100011;
#10000;
	data_in <= 24'b010111110101000001001101;
#10000;
	data_in <= 24'b000010110000100000000000;
#10000;
	data_in <= 24'b000011010000100100001000;
#10000;
	data_in <= 24'b000010000000010100001110;
#10000;
	data_in <= 24'b000001110000011100010101;
#10000;
	data_in <= 24'b000001100000101100011010;
#10000;
	data_in <= 24'b000010110000111100011010;
#10000;
	data_in <= 24'b001010010010100000101010;
#10000;
	data_in <= 24'b011111010111000101101011;
#10000;
	data_in <= 24'b000011110000110100000101;
#10000;
	data_in <= 24'b000100000000111100001011;
#10000;
	data_in <= 24'b000010000000100100001101;
#10000;
	data_in <= 24'b000001010000011100010001;
#10000;
	data_in <= 24'b000011010001001100100000;
#10000;
	data_in <= 24'b000100010001011000011111;
#10000;
	data_in <= 24'b001000100010010000100100;
#10000;
	data_in <= 24'b010011100100011100111110;
#10000;
	data_in <= 24'b000001010000100100001010;
#10000;
	data_in <= 24'b000001000000100000001001;
#10000;
	data_in <= 24'b000010100000111000001111;
#10000;
	data_in <= 24'b000101010001100100011110;
#10000;
	data_in <= 24'b000110110001111100101010;
#10000;
	data_in <= 24'b000010010000101100010101;
#10000;
	data_in <= 24'b000110100001101100011001;
#10000;
	data_in <= 24'b001101000011001000101000;
#10000;
	data_in <= 24'b001001100010111000111011;
#10000;
	data_in <= 24'b001010110011010000111110;
#10000;
	data_in <= 24'b001101010011110101000100;
#10000;
	data_in <= 24'b001110110100001001001011;
#10000;
	data_in <= 24'b010010000100110101011100;
#10000;
	data_in <= 24'b010000100100010101010100;
#10000;
	data_in <= 24'b010110100101110101100101;
#10000;
	data_in <= 24'b010111010110000001100100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001011100001111000001101;
#10000;
	data_in <= 24'b001110100010110000010110;
#10000;
	data_in <= 24'b001110000010111000010110;
#10000;
	data_in <= 24'b001010100010010000010001;
#10000;
	data_in <= 24'b001000100001110100011010;
#10000;
	data_in <= 24'b001010010010010000100101;
#10000;
	data_in <= 24'b001100000010101000100011;
#10000;
	data_in <= 24'b001101000011000100101001;
#10000;
	data_in <= 24'b100100100111110001101010;
#10000;
	data_in <= 24'b100101000111111101100000;
#10000;
	data_in <= 24'b100110111000110101100011;
#10000;
	data_in <= 24'b010000010011011100010101;
#10000;
	data_in <= 24'b001010000001111000010111;
#10000;
	data_in <= 24'b001000010001011100010111;
#10000;
	data_in <= 24'b001101110010111000100100;
#10000;
	data_in <= 24'b000110010001011000001000;
#10000;
	data_in <= 24'b111011101101001011000001;
#10000;
	data_in <= 24'b110100111011001110001111;
#10000;
	data_in <= 24'b110001111010111101110011;
#10000;
	data_in <= 24'b100011110111101001000011;
#10000;
	data_in <= 24'b001011100001010000000110;
#10000;
	data_in <= 24'b011011100101011101010101;
#10000;
	data_in <= 24'b101100101010001010010001;
#10000;
	data_in <= 24'b000111100001100000000001;
#10000;
	data_in <= 24'b100000100110010001010011;
#10000;
	data_in <= 24'b100110000111010001001110;
#10000;
	data_in <= 24'b101110001001110001010101;
#10000;
	data_in <= 24'b101010111001000101001111;
#10000;
	data_in <= 24'b010000100010001000001111;
#10000;
	data_in <= 24'b100001110110110001101000;
#10000;
	data_in <= 24'b011011000101101101000110;
#10000;
	data_in <= 24'b001010100010001100001010;
#10000;
	data_in <= 24'b100001010110101101011011;
#10000;
	data_in <= 24'b101000001000000101011010;
#10000;
	data_in <= 24'b101111011010011001011010;
#10000;
	data_in <= 24'b100110101000001100111111;
#10000;
	data_in <= 24'b010101100011101100100111;
#10000;
	data_in <= 24'b010101010011111000111100;
#10000;
	data_in <= 24'b001111100011010100100001;
#10000;
	data_in <= 24'b001101000011000000011000;
#10000;
	data_in <= 24'b100001010111000001100001;
#10000;
	data_in <= 24'b101000111000101001101000;
#10000;
	data_in <= 24'b101101001010001101100000;
#10000;
	data_in <= 24'b100111011000111001010000;
#10000;
	data_in <= 24'b001111000010100000010110;
#10000;
	data_in <= 24'b001100110010001000011111;
#10000;
	data_in <= 24'b001100010010110100011010;
#10000;
	data_in <= 24'b001011000010100100010100;
#10000;
	data_in <= 24'b010100110100011100111011;
#10000;
	data_in <= 24'b001110100010110100010011;
#10000;
	data_in <= 24'b101000011001100101101010;
#10000;
	data_in <= 24'b100011001000011001011001;
#10000;
	data_in <= 24'b011001110101110001001110;
#10000;
	data_in <= 24'b011101100110111001100111;
#10000;
	data_in <= 24'b011010010110100101010111;
#10000;
	data_in <= 24'b011011110111000101011011;
#10000;
	data_in <= 24'b011100100111010001110101;
#10000;
	data_in <= 24'b100010101000101110000111;
#10000;
	data_in <= 24'b100100111001101010001011;
#10000;
	data_in <= 24'b100101001001110010010001;
#10000;
	data_in <= 24'b100110001001110110100000;
#10000;
	data_in <= 24'b101100001011010110111110;
#10000;
	data_in <= 24'b101101101100000011000000;
#10000;
	data_in <= 24'b101100101100000010111110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001000100010001100011111;
#10000;
	data_in <= 24'b001000010010001100100100;
#10000;
	data_in <= 24'b001001010010000100100111;
#10000;
	data_in <= 24'b000110110001010000011011;
#10000;
	data_in <= 24'b000111100001100000011001;
#10000;
	data_in <= 24'b000111000001010100010010;
#10000;
	data_in <= 24'b000110000001000000010000;
#10000;
	data_in <= 24'b000100110000111000001101;
#10000;
	data_in <= 24'b000011010001000000000111;
#10000;
	data_in <= 24'b000010010000111000001100;
#10000;
	data_in <= 24'b000010110000011100001100;
#10000;
	data_in <= 24'b000011100000100100001011;
#10000;
	data_in <= 24'b000111100001011100010100;
#10000;
	data_in <= 24'b000101110001000100001100;
#10000;
	data_in <= 24'b000101100000111100001100;
#10000;
	data_in <= 24'b000100010000110100001100;
#10000;
	data_in <= 24'b000110000001101100001011;
#10000;
	data_in <= 24'b000111010010010000010111;
#10000;
	data_in <= 24'b000110000001100000001100;
#10000;
	data_in <= 24'b010000010011111100110100;
#10000;
	data_in <= 24'b010001000011111000110011;
#10000;
	data_in <= 24'b001011000010010100011100;
#10000;
	data_in <= 24'b000110100001000100001101;
#10000;
	data_in <= 24'b000110100001010100010100;
#10000;
	data_in <= 24'b001011000010101000011000;
#10000;
	data_in <= 24'b001010100010100100011011;
#10000;
	data_in <= 24'b001101000011001000100000;
#10000;
	data_in <= 24'b011100010110110101011011;
#10000;
	data_in <= 24'b010001110100000100110110;
#10000;
	data_in <= 24'b001011100010100000100001;
#10000;
	data_in <= 24'b000110100001010100010100;
#10000;
	data_in <= 24'b001000000001110100011111;
#10000;
	data_in <= 24'b001110100010111000100100;
#10000;
	data_in <= 24'b001011110010001000011010;
#10000;
	data_in <= 24'b011111010111001101100010;
#10000;
	data_in <= 24'b100100011000100001111010;
#10000;
	data_in <= 24'b010101100100110101001001;
#10000;
	data_in <= 24'b010010110100011001001000;
#10000;
	data_in <= 24'b001111110011111001000111;
#10000;
	data_in <= 24'b001100000011011001000011;
#10000;
	data_in <= 24'b001101100010110000100010;
#10000;
	data_in <= 24'b001000010001010000001100;
#10000;
	data_in <= 24'b101011111010010110010100;
#10000;
	data_in <= 24'b100100101000101101111100;
#10000;
	data_in <= 24'b010110110101010001010001;
#10000;
	data_in <= 24'b011000000101111001100100;
#10000;
	data_in <= 24'b011001000110100001110011;
#10000;
	data_in <= 24'b001011110011100101001011;
#10000;
	data_in <= 24'b011010100110011101011000;
#10000;
	data_in <= 24'b011101110111010001100101;
#10000;
	data_in <= 24'b101000111010001010001110;
#10000;
	data_in <= 24'b011010000110100001011000;
#10000;
	data_in <= 24'b010101100101001101001110;
#10000;
	data_in <= 24'b001111110100000001000100;
#10000;
	data_in <= 24'b001001100010101000110101;
#10000;
	data_in <= 24'b000111000010001100110110;
#10000;
	data_in <= 24'b101110101100101011001001;
#10000;
	data_in <= 24'b101110011100101111001010;
#10000;
	data_in <= 24'b100100111010010110100100;
#10000;
	data_in <= 24'b100010001001101110011110;
#10000;
	data_in <= 24'b010110010110110001110100;
#10000;
	data_in <= 24'b010000100101011001100111;
#10000;
	data_in <= 24'b001111000101001101101001;
#10000;
	data_in <= 24'b001101110101001001101100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000101000001001000010010;
#10000;
	data_in <= 24'b001001100010001100100101;
#10000;
	data_in <= 24'b001110100011100100111011;
#10000;
	data_in <= 24'b001101110011001100111000;
#10000;
	data_in <= 24'b001110010011000100111000;
#10000;
	data_in <= 24'b001101110010110000101111;
#10000;
	data_in <= 24'b001011110010001100011111;
#10000;
	data_in <= 24'b001100100010011000011100;
#10000;
	data_in <= 24'b000011110000110000001110;
#10000;
	data_in <= 24'b000001010000010100001011;
#10000;
	data_in <= 24'b000001110000101000001111;
#10000;
	data_in <= 24'b000100100001000100011010;
#10000;
	data_in <= 24'b000110100001010000011111;
#10000;
	data_in <= 24'b000100010000100100010000;
#10000;
	data_in <= 24'b000111000001000000010000;
#10000;
	data_in <= 24'b000101010000100100000101;
#10000;
	data_in <= 24'b000100000000101100001101;
#10000;
	data_in <= 24'b000011100000110000010010;
#10000;
	data_in <= 24'b000101010001010000011110;
#10000;
	data_in <= 24'b000111110001111000101000;
#10000;
	data_in <= 24'b001000000001110000100111;
#10000;
	data_in <= 24'b001010010010000100101011;
#10000;
	data_in <= 24'b000110000000111000010100;
#10000;
	data_in <= 24'b001111010010110100111000;
#10000;
	data_in <= 24'b000101000001011000011110;
#10000;
	data_in <= 24'b000010110000111000011100;
#10000;
	data_in <= 24'b000010000000110100011100;
#10000;
	data_in <= 24'b000001010000101000011001;
#10000;
	data_in <= 24'b000000010000010000010010;
#10000;
	data_in <= 24'b000011010000110100011001;
#10000;
	data_in <= 24'b001001110010001000110001;
#10000;
	data_in <= 24'b011111010111001110001010;
#10000;
	data_in <= 24'b010010000101010001100110;
#10000;
	data_in <= 24'b100001101001011010101101;
#10000;
	data_in <= 24'b100101001010010110111111;
#10000;
	data_in <= 24'b100111001010101111000101;
#10000;
	data_in <= 24'b100101001010001110110110;
#10000;
	data_in <= 24'b000101100010000100110101;
#10000;
	data_in <= 24'b001001010010100101000101;
#10000;
	data_in <= 24'b010011010101001001110011;
#10000;
	data_in <= 24'b001001100011011001001101;
#10000;
	data_in <= 24'b011111011001001010101110;
#10000;
	data_in <= 24'b100011101010001111000010;
#10000;
	data_in <= 24'b100001101001111010111010;
#10000;
	data_in <= 24'b011010101000000010011001;
#10000;
	data_in <= 24'b000000000000111000100111;
#10000;
	data_in <= 24'b010000110100111101110001;
#10000;
	data_in <= 24'b011000100111010010011001;
#10000;
	data_in <= 24'b001000100011000001000111;
#10000;
	data_in <= 24'b000100010010010000111111;
#10000;
	data_in <= 24'b000001100001101100111010;
#10000;
	data_in <= 24'b000000000001010000110010;
#10000;
	data_in <= 24'b000000000000001100011101;
#10000;
	data_in <= 24'b000000000001001100101101;
#10000;
	data_in <= 24'b010101110110110110010000;
#10000;
	data_in <= 24'b010101100111010010010111;
#10000;
	data_in <= 24'b001110110101100101110110;
#10000;
	data_in <= 24'b001101110101100101110111;
#10000;
	data_in <= 24'b010011000111001010010010;
#10000;
	data_in <= 24'b010011010111001110010011;
#10000;
	data_in <= 24'b010101000111101010011000;
#10000;
	data_in <= 24'b010011100111010010010010;
#10000;
	data_in <= 24'b011011001000111110110000;
#10000;
	data_in <= 24'b011100011001100010111000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001101010010011100011011;
#10000;
	data_in <= 24'b001100110010011100011101;
#10000;
	data_in <= 24'b001100100010100000100001;
#10000;
	data_in <= 24'b001101100010101000100100;
#10000;
	data_in <= 24'b010011010011101000101101;
#10000;
	data_in <= 24'b010100000011010100100111;
#10000;
	data_in <= 24'b011000010011111000110001;
#10000;
	data_in <= 24'b011011000100011001000001;
#10000;
	data_in <= 24'b001001010001011000010100;
#10000;
	data_in <= 24'b010000110011001100110100;
#10000;
	data_in <= 24'b010000100011010000110110;
#10000;
	data_in <= 24'b010001100011001100110000;
#10000;
	data_in <= 24'b010010110011001000100010;
#10000;
	data_in <= 24'b010101100011011000011111;
#10000;
	data_in <= 24'b011000100011100100100011;
#10000;
	data_in <= 24'b011011010100000100110100;
#10000;
	data_in <= 24'b011100000101100001110000;
#10000;
	data_in <= 24'b010011010011000001001010;
#10000;
	data_in <= 24'b010010010010100000111101;
#10000;
	data_in <= 24'b010101000010111000110100;
#10000;
	data_in <= 24'b011011000100000000101111;
#10000;
	data_in <= 24'b011011110100000000100001;
#10000;
	data_in <= 24'b011011110011111100011101;
#10000;
	data_in <= 24'b011001000011011100011100;
#10000;
	data_in <= 24'b100011010111111110100011;
#10000;
	data_in <= 24'b011100110101110010000010;
#10000;
	data_in <= 24'b011111100101110101111000;
#10000;
	data_in <= 24'b100011110110010001101101;
#10000;
	data_in <= 24'b100011110101101101001010;
#10000;
	data_in <= 24'b110101011001111101111110;
#10000;
	data_in <= 24'b110000001000111101100111;
#10000;
	data_in <= 24'b011011100100010100100101;
#10000;
	data_in <= 24'b011111101000101010101110;
#10000;
	data_in <= 24'b100111111010010011000101;
#10000;
	data_in <= 24'b101100111010001110111011;
#10000;
	data_in <= 24'b101010111000101010010001;
#10000;
	data_in <= 24'b101000110111010101100011;
#10000;
	data_in <= 24'b111111111101010110110101;
#10000;
	data_in <= 24'b111111111101111110111010;
#10000;
	data_in <= 24'b101011001000110001101111;
#10000;
	data_in <= 24'b100011001010101011001101;
#10000;
	data_in <= 24'b101000001011011111010111;
#10000;
	data_in <= 24'b011111100111101110010101;
#10000;
	data_in <= 24'b100101000111110110001011;
#10000;
	data_in <= 24'b011000100011101000110101;
#10000;
	data_in <= 24'b101111101001001110000000;
#10000;
	data_in <= 24'b111000001011111010100111;
#10000;
	data_in <= 24'b111111001110010111010110;
#10000;
	data_in <= 24'b100101101100000011100011;
#10000;
	data_in <= 24'b100110011011111011100000;
#10000;
	data_in <= 24'b010111010110010110001010;
#10000;
	data_in <= 24'b010100010100001001100001;
#10000;
	data_in <= 24'b011011010100110101011110;
#10000;
	data_in <= 24'b101010111000011010010000;
#10000;
	data_in <= 24'b101000101000100010001110;
#10000;
	data_in <= 24'b111111111111101111111111;
#10000;
	data_in <= 24'b011010001001101010111000;
#10000;
	data_in <= 24'b011011101001101010111001;
#10000;
	data_in <= 24'b100101001010011111001010;
#10000;
	data_in <= 24'b010111010101110001111110;
#10000;
	data_in <= 24'b010001110011010001001111;
#10000;
	data_in <= 24'b100101100111111010010110;
#10000;
	data_in <= 24'b100010010111110110001111;
#10000;
	data_in <= 24'b110101111101011111101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011010100011001001110;
#10000;
	data_in <= 24'b011010110100011101010111;
#10000;
	data_in <= 24'b011011100101000101100000;
#10000;
	data_in <= 24'b011010100101001001011110;
#10000;
	data_in <= 24'b011011010101011101011100;
#10000;
	data_in <= 24'b011011100101101001011111;
#10000;
	data_in <= 24'b011010000101001001011110;
#10000;
	data_in <= 24'b011001000101001101100000;
#10000;
	data_in <= 24'b011101110100111001010101;
#10000;
	data_in <= 24'b011110100101011001100110;
#10000;
	data_in <= 24'b011100000101010001100111;
#10000;
	data_in <= 24'b011011100101100101101000;
#10000;
	data_in <= 24'b011101100110010001101011;
#10000;
	data_in <= 24'b011101000110010001101011;
#10000;
	data_in <= 24'b011011000101110101101011;
#10000;
	data_in <= 24'b010111110101011101101000;
#10000;
	data_in <= 24'b011001000011111000111010;
#10000;
	data_in <= 24'b011010110100110001010101;
#10000;
	data_in <= 24'b011001010100101101011011;
#10000;
	data_in <= 24'b011010100101010001100110;
#10000;
	data_in <= 24'b011010110101100101100110;
#10000;
	data_in <= 24'b011100100110010001110000;
#10000;
	data_in <= 24'b011011110110010101110110;
#10000;
	data_in <= 24'b100110101001110010101110;
#10000;
	data_in <= 24'b010111110100000000110111;
#10000;
	data_in <= 24'b010100000011100001000000;
#10000;
	data_in <= 24'b010111010100010001011000;
#10000;
	data_in <= 24'b100011100111100110001111;
#10000;
	data_in <= 24'b100110111000100110011010;
#10000;
	data_in <= 24'b110010011011110011001100;
#10000;
	data_in <= 24'b101111101011101011001101;
#10000;
	data_in <= 24'b110010111101001011100101;
#10000;
	data_in <= 24'b100100000111101001110101;
#10000;
	data_in <= 24'b010010100011100101000110;
#10000;
	data_in <= 24'b100010110111011010001111;
#10000;
	data_in <= 24'b111001011101001011101101;
#10000;
	data_in <= 24'b101111001010100110111110;
#10000;
	data_in <= 24'b101111001011000011000010;
#10000;
	data_in <= 24'b110011011100101111011111;
#10000;
	data_in <= 24'b110011001101010111101001;
#10000;
	data_in <= 24'b110010001011110011000010;
#10000;
	data_in <= 24'b010101010100111101100010;
#10000;
	data_in <= 24'b101010101010000110111100;
#10000;
	data_in <= 24'b111001011101100111110101;
#10000;
	data_in <= 24'b110010011011110111010011;
#10000;
	data_in <= 24'b110001101100000011010001;
#10000;
	data_in <= 24'b110001001100100011011010;
#10000;
	data_in <= 24'b110001111101011011101001;
#10000;
	data_in <= 24'b110010001100100111011101;
#10000;
	data_in <= 24'b011100110111101010010011;
#10000;
	data_in <= 24'b110000101100011011100010;
#10000;
	data_in <= 24'b111000001110010011111100;
#10000;
	data_in <= 24'b110110111101111011101101;
#10000;
	data_in <= 24'b101111101100100011010010;
#10000;
	data_in <= 24'b101001111011110011000100;
#10000;
	data_in <= 24'b111000111111110111111111;
#10000;
	data_in <= 24'b110011001101101011110001;
#10000;
	data_in <= 24'b100111011011001111001100;
#10000;
	data_in <= 24'b101100101100010011011011;
#10000;
	data_in <= 24'b110110101110101111111110;
#10000;
	data_in <= 24'b111011011111110111111111;
#10000;
	data_in <= 24'b110101101110101011110101;
#10000;
	data_in <= 24'b101101101101010111011110;
#10000;
	data_in <= 24'b110100001111000111111111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011011010110011101110010;
#10000;
	data_in <= 24'b010111010101011001011101;
#10000;
	data_in <= 24'b011011000101011001011011;
#10000;
	data_in <= 24'b011101110101011001011010;
#10000;
	data_in <= 24'b100000010101101001011000;
#10000;
	data_in <= 24'b011111100101100101010001;
#10000;
	data_in <= 24'b100000100110000001010011;
#10000;
	data_in <= 24'b011111100110000001001111;
#10000;
	data_in <= 24'b110101011101110011101011;
#10000;
	data_in <= 24'b100101101001100110100111;
#10000;
	data_in <= 24'b011000010101000001011101;
#10000;
	data_in <= 24'b100000000110001101101100;
#10000;
	data_in <= 24'b100010110110011101101101;
#10000;
	data_in <= 24'b100011000110101001101011;
#10000;
	data_in <= 24'b100001000110101101100111;
#10000;
	data_in <= 24'b100001000110111101100111;
#10000;
	data_in <= 24'b101110111100101111011011;
#10000;
	data_in <= 24'b101001011011010011000100;
#10000;
	data_in <= 24'b001110010011001001000001;
#10000;
	data_in <= 24'b010001000010111100111110;
#10000;
	data_in <= 24'b010010010011000100111101;
#10000;
	data_in <= 24'b001110110010100000110001;
#10000;
	data_in <= 24'b001011110010010000101100;
#10000;
	data_in <= 24'b000111010001100100011110;
#10000;
	data_in <= 24'b111001101111110011111111;
#10000;
	data_in <= 24'b100101011010100110111011;
#10000;
	data_in <= 24'b001010000010011000111010;
#10000;
	data_in <= 24'b001100010010010100111001;
#10000;
	data_in <= 24'b001010110001110100101111;
#10000;
	data_in <= 24'b000111000001010000100101;
#10000;
	data_in <= 24'b000101010001101000101001;
#10000;
	data_in <= 24'b000101000001110100101011;
#10000;
	data_in <= 24'b110111111111011011111111;
#10000;
	data_in <= 24'b100000101001011010101111;
#10000;
	data_in <= 24'b001011100010110101000111;
#10000;
	data_in <= 24'b001100000010011101000001;
#10000;
	data_in <= 24'b001000000001101000110011;
#10000;
	data_in <= 24'b000100000001001100101000;
#10000;
	data_in <= 24'b000111000010110101000000;
#10000;
	data_in <= 24'b010010010101111101110001;
#10000;
	data_in <= 24'b101011111100010011011111;
#10000;
	data_in <= 24'b001111100101000001101101;
#10000;
	data_in <= 24'b001011010010111101001101;
#10000;
	data_in <= 24'b001001110010001101000000;
#10000;
	data_in <= 24'b001011000010110101001001;
#10000;
	data_in <= 24'b011111111000101110100011;
#10000;
	data_in <= 24'b011100001000100010011110;
#10000;
	data_in <= 24'b010000100110001001110101;
#10000;
	data_in <= 24'b100110111011000011001011;
#10000;
	data_in <= 24'b001101110100010001100100;
#10000;
	data_in <= 24'b010101100101100101111000;
#10000;
	data_in <= 24'b010001100100100001100110;
#10000;
	data_in <= 24'b100011011001001110110000;
#10000;
	data_in <= 24'b101111011100111011101000;
#10000;
	data_in <= 24'b011100101001000110100110;
#10000;
	data_in <= 24'b101110101101101111101111;
#10000;
	data_in <= 24'b101000111100000111011100;
#10000;
	data_in <= 24'b011100001000100110101001;
#10000;
	data_in <= 24'b101000011011010111010100;
#10000;
	data_in <= 24'b100000111001011110110110;
#10000;
	data_in <= 24'b101011001100011011100100;
#10000;
	data_in <= 24'b110000101110010111111111;
#10000;
	data_in <= 24'b101011011101100111110001;
#10000;
	data_in <= 24'b101100011101110111110101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100000000110001001001111;
#10000;
	data_in <= 24'b100001100110101001010010;
#10000;
	data_in <= 24'b100010010110111001010100;
#10000;
	data_in <= 24'b100010010110110101001111;
#10000;
	data_in <= 24'b100011100111001001010011;
#10000;
	data_in <= 24'b100011110111000001001111;
#10000;
	data_in <= 24'b100101110111010001010010;
#10000;
	data_in <= 24'b100110100111010001010001;
#10000;
	data_in <= 24'b011110110110100101011110;
#10000;
	data_in <= 24'b011000100100111101000010;
#10000;
	data_in <= 24'b011000100100111101000000;
#10000;
	data_in <= 24'b010111010100100100111000;
#10000;
	data_in <= 24'b010111110100100100110111;
#10000;
	data_in <= 24'b011001010100110100111001;
#10000;
	data_in <= 24'b011100000101001100111110;
#10000;
	data_in <= 24'b011111110110000101001000;
#10000;
	data_in <= 24'b000111100001100000011101;
#10000;
	data_in <= 24'b011001110110000001100101;
#10000;
	data_in <= 24'b001000010001010100011011;
#10000;
	data_in <= 24'b000100110000010100001011;
#10000;
	data_in <= 24'b000101100000011100001011;
#10000;
	data_in <= 24'b000100100000010000000110;
#10000;
	data_in <= 24'b000110010000100000001011;
#10000;
	data_in <= 24'b000110010000101000001000;
#10000;
	data_in <= 24'b001111100100010101010100;
#10000;
	data_in <= 24'b010111000101111101101110;
#10000;
	data_in <= 24'b000111110001100100101100;
#10000;
	data_in <= 24'b000110010000111100100000;
#10000;
	data_in <= 24'b000110000000111000011111;
#10000;
	data_in <= 24'b000110100001000000100000;
#10000;
	data_in <= 24'b000100100000101100011000;
#10000;
	data_in <= 24'b000100010000110100011000;
#10000;
	data_in <= 24'b001001000011100001001010;
#10000;
	data_in <= 24'b000100010001110000110000;
#10000;
	data_in <= 24'b001101010011011001001010;
#10000;
	data_in <= 24'b000101110001001000100111;
#10000;
	data_in <= 24'b000010110000100000011000;
#10000;
	data_in <= 24'b000011000000110000011010;
#10000;
	data_in <= 24'b000011010001000100011100;
#10000;
	data_in <= 24'b000010000000111000011001;
#10000;
	data_in <= 24'b000111000011010101001001;
#10000;
	data_in <= 24'b000010110001110000110001;
#10000;
	data_in <= 24'b001111110100001001010111;
#10000;
	data_in <= 24'b000111110001110100110000;
#10000;
	data_in <= 24'b000101000001001100100011;
#10000;
	data_in <= 24'b000011110001001100011110;
#10000;
	data_in <= 24'b000100010001101000100011;
#10000;
	data_in <= 24'b000001100001000100011001;
#10000;
	data_in <= 24'b011001111000000010010100;
#10000;
	data_in <= 24'b000000000000110100100000;
#10000;
	data_in <= 24'b000100010001011100101010;
#10000;
	data_in <= 24'b000111010001110100101101;
#10000;
	data_in <= 24'b000110010001101100100101;
#10000;
	data_in <= 24'b000110010001111100100100;
#10000;
	data_in <= 24'b000010010001010100010111;
#10000;
	data_in <= 24'b000100100001101100011110;
#10000;
	data_in <= 24'b010001110110100010000010;
#10000;
	data_in <= 24'b000000000000100000100010;
#10000;
	data_in <= 24'b000011100001110100110111;
#10000;
	data_in <= 24'b000011110001110000110010;
#10000;
	data_in <= 24'b000011000001100000101010;
#10000;
	data_in <= 24'b000000110001001100100000;
#10000;
	data_in <= 24'b000000000000111100011000;
#10000;
	data_in <= 24'b000001100001010000100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100110010111001001001011;
#10000;
	data_in <= 24'b100110110111001101001001;
#10000;
	data_in <= 24'b100110010111000001001001;
#10000;
	data_in <= 24'b100110010110111101000101;
#10000;
	data_in <= 24'b100110100110111001000101;
#10000;
	data_in <= 24'b100110010110111001000011;
#10000;
	data_in <= 24'b100101100110100100111110;
#10000;
	data_in <= 24'b100100000110001000111001;
#10000;
	data_in <= 24'b100001000110011001001001;
#10000;
	data_in <= 24'b100100110111010001010101;
#10000;
	data_in <= 24'b101000111000000101100011;
#10000;
	data_in <= 24'b101010011000100001100111;
#10000;
	data_in <= 24'b101010111000011001100100;
#10000;
	data_in <= 24'b101001000111111101011101;
#10000;
	data_in <= 24'b100111010111011101010101;
#10000;
	data_in <= 24'b100101110111000101001111;
#10000;
	data_in <= 24'b000111000000111100000111;
#10000;
	data_in <= 24'b001001100001100000001100;
#10000;
	data_in <= 24'b001110000010100000011100;
#10000;
	data_in <= 24'b010011110011111100110010;
#10000;
	data_in <= 24'b011010110101100001001001;
#10000;
	data_in <= 24'b100000000110111001011101;
#10000;
	data_in <= 24'b100011010111100101100111;
#10000;
	data_in <= 24'b100100100111110101101000;
#10000;
	data_in <= 24'b000100000000111000010100;
#10000;
	data_in <= 24'b000011010000110000001110;
#10000;
	data_in <= 24'b000010010000011000001000;
#10000;
	data_in <= 24'b000001010000000000000001;
#10000;
	data_in <= 24'b000001110000001000000000;
#10000;
	data_in <= 24'b000100110000110100001000;
#10000;
	data_in <= 24'b001000110001101100010100;
#10000;
	data_in <= 24'b001100000010011100011110;
#10000;
	data_in <= 24'b000010000000110000010111;
#10000;
	data_in <= 24'b000010110000111100011010;
#10000;
	data_in <= 24'b000011110001000100011011;
#10000;
	data_in <= 24'b000100000001001000011010;
#10000;
	data_in <= 24'b000011100000111000010100;
#10000;
	data_in <= 24'b000011000000101100001111;
#10000;
	data_in <= 24'b000010110000101100001011;
#10000;
	data_in <= 24'b000011100000110000001011;
#10000;
	data_in <= 24'b000010010000111100011100;
#10000;
	data_in <= 24'b000001100000100100010111;
#10000;
	data_in <= 24'b000001010000011100010010;
#10000;
	data_in <= 24'b000001110000100100010100;
#10000;
	data_in <= 24'b000010110000110000010110;
#10000;
	data_in <= 24'b000011000000111000010110;
#10000;
	data_in <= 24'b000011010000110100010011;
#10000;
	data_in <= 24'b000010110000110000010000;
#10000;
	data_in <= 24'b000111110010000100101001;
#10000;
	data_in <= 24'b001001000010001100101100;
#10000;
	data_in <= 24'b001010100010011100110000;
#10000;
	data_in <= 24'b001010010010011000101111;
#10000;
	data_in <= 24'b001001010010000100100111;
#10000;
	data_in <= 24'b000111100001101000100000;
#10000;
	data_in <= 24'b000110100001011000011011;
#10000;
	data_in <= 24'b000110110001011100011100;
#10000;
	data_in <= 24'b000111000010010100110011;
#10000;
	data_in <= 24'b000101110001101100101101;
#10000;
	data_in <= 24'b000100000001010000100110;
#10000;
	data_in <= 24'b000011010001000100100011;
#10000;
	data_in <= 24'b000011100001000100100000;
#10000;
	data_in <= 24'b000011010001000000011111;
#10000;
	data_in <= 24'b000011010001000000011111;
#10000;
	data_in <= 24'b000011010001000000011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100011000101111100111001;
#10000;
	data_in <= 24'b100010000101101100110110;
#10000;
	data_in <= 24'b100000100101010100110011;
#10000;
	data_in <= 24'b011111010101001000110001;
#10000;
	data_in <= 24'b011101110100110100110000;
#10000;
	data_in <= 24'b011100000100100000101100;
#10000;
	data_in <= 24'b011010100100001000101001;
#10000;
	data_in <= 24'b011010000100000100100101;
#10000;
	data_in <= 24'b100010100110010001000010;
#10000;
	data_in <= 24'b100001100110000001000000;
#10000;
	data_in <= 24'b100000000101101100111111;
#10000;
	data_in <= 24'b011110110101011000111100;
#10000;
	data_in <= 24'b011100110100111100110111;
#10000;
	data_in <= 24'b011011000100101000110011;
#10000;
	data_in <= 24'b011010000100011100110011;
#10000;
	data_in <= 24'b011010000100100100110100;
#10000;
	data_in <= 24'b100011100111100101100100;
#10000;
	data_in <= 24'b100000010110101101011001;
#10000;
	data_in <= 24'b011011100101101001001000;
#10000;
	data_in <= 24'b011000010100110100111100;
#10000;
	data_in <= 24'b010101100100001100110100;
#10000;
	data_in <= 24'b010011000011101100101110;
#10000;
	data_in <= 24'b010001100011010100101000;
#10000;
	data_in <= 24'b010000100011000000100101;
#10000;
	data_in <= 24'b010010100100000100111000;
#10000;
	data_in <= 24'b001110000010111100100101;
#10000;
	data_in <= 24'b001000010001100000001111;
#10000;
	data_in <= 24'b000100010000101000000001;
#10000;
	data_in <= 24'b000011010000010100000000;
#10000;
	data_in <= 24'b000011010000011100000000;
#10000;
	data_in <= 24'b000011110000100100000010;
#10000;
	data_in <= 24'b000100000000101000000101;
#10000;
	data_in <= 24'b000001100000010000000011;
#10000;
	data_in <= 24'b000010010000011100000110;
#10000;
	data_in <= 24'b000011100000110000001011;
#10000;
	data_in <= 24'b000011110001000000001110;
#10000;
	data_in <= 24'b000100000001000100001111;
#10000;
	data_in <= 24'b000010110000111000001100;
#10000;
	data_in <= 24'b000010010000110000001010;
#10000;
	data_in <= 24'b000001110000110000001011;
#10000;
	data_in <= 24'b000011110001000100010010;
#10000;
	data_in <= 24'b000011100001000000010001;
#10000;
	data_in <= 24'b000011100001000000010001;
#10000;
	data_in <= 24'b000011000001000000010001;
#10000;
	data_in <= 24'b000010110000111100010000;
#10000;
	data_in <= 24'b000010010000111000010001;
#10000;
	data_in <= 24'b000010100000111100010010;
#10000;
	data_in <= 24'b000010100001000100010100;
#10000;
	data_in <= 24'b000111100001101000011111;
#10000;
	data_in <= 24'b000101110001011000011010;
#10000;
	data_in <= 24'b000101000001001100010111;
#10000;
	data_in <= 24'b000100100001001100010111;
#10000;
	data_in <= 24'b000100110001010000011000;
#10000;
	data_in <= 24'b000011110001001000010111;
#10000;
	data_in <= 24'b000011010001000000010101;
#10000;
	data_in <= 24'b000010110000110100010101;
#10000;
	data_in <= 24'b000010010000111000011101;
#10000;
	data_in <= 24'b000010110001000000011111;
#10000;
	data_in <= 24'b000011100001001100100010;
#10000;
	data_in <= 24'b000100100001011100100110;
#10000;
	data_in <= 24'b000100010001100000101001;
#10000;
	data_in <= 24'b000100000001011100101000;
#10000;
	data_in <= 24'b000100000001100000101001;
#10000;
	data_in <= 24'b000100110001101000101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011001110100001100100101;
#10000;
	data_in <= 24'b011000110100000000011111;
#10000;
	data_in <= 24'b010111110011111000011101;
#10000;
	data_in <= 24'b011000000011111100011110;
#10000;
	data_in <= 24'b011000010011111100100001;
#10000;
	data_in <= 24'b010111110011111100100010;
#10000;
	data_in <= 24'b011000010100000000100110;
#10000;
	data_in <= 24'b011000010100001100101000;
#10000;
	data_in <= 24'b011000010100000100101010;
#10000;
	data_in <= 24'b011000010100001000101011;
#10000;
	data_in <= 24'b011000100100001100101100;
#10000;
	data_in <= 24'b011000010100010100101101;
#10000;
	data_in <= 24'b010111100100001000101010;
#10000;
	data_in <= 24'b010110010011111000101001;
#10000;
	data_in <= 24'b010101110011110000101000;
#10000;
	data_in <= 24'b010101000011110000101010;
#10000;
	data_in <= 24'b010011100011100100110001;
#10000;
	data_in <= 24'b010011110011100100110011;
#10000;
	data_in <= 24'b010011000011011000110000;
#10000;
	data_in <= 24'b010000000010110100100110;
#10000;
	data_in <= 24'b001100110010000000011001;
#10000;
	data_in <= 24'b001001100001001100001110;
#10000;
	data_in <= 24'b000111000000110000000110;
#10000;
	data_in <= 24'b000101100000011100000100;
#10000;
	data_in <= 24'b000100110000100100001001;
#10000;
	data_in <= 24'b000101110000110000001110;
#10000;
	data_in <= 24'b000110000000110100001111;
#10000;
	data_in <= 24'b000100110000100000001010;
#10000;
	data_in <= 24'b000011110000010000000110;
#10000;
	data_in <= 24'b000011000000010000000101;
#10000;
	data_in <= 24'b000011000000001100000110;
#10000;
	data_in <= 24'b000010100000001100000110;
#10000;
	data_in <= 24'b000001100000100000001000;
#10000;
	data_in <= 24'b000010000000101000001010;
#10000;
	data_in <= 24'b000001110000100100001001;
#10000;
	data_in <= 24'b000001000000011000000110;
#10000;
	data_in <= 24'b000001000000011000000110;
#10000;
	data_in <= 24'b000010010000100100001001;
#10000;
	data_in <= 24'b000010110000101100001011;
#10000;
	data_in <= 24'b000010110000101100001011;
#10000;
	data_in <= 24'b000001110000111000010001;
#10000;
	data_in <= 24'b000001110000111000010001;
#10000;
	data_in <= 24'b000010000000110100010000;
#10000;
	data_in <= 24'b000001110000110000001111;
#10000;
	data_in <= 24'b000010000000110100010000;
#10000;
	data_in <= 24'b000010010000111000001111;
#10000;
	data_in <= 24'b000010100000111000001111;
#10000;
	data_in <= 24'b000010000000110000001101;
#10000;
	data_in <= 24'b000011100000111100011001;
#10000;
	data_in <= 24'b000011010000111000011000;
#10000;
	data_in <= 24'b000011010000111000011000;
#10000;
	data_in <= 24'b000011110001000000011010;
#10000;
	data_in <= 24'b000011110001000000011010;
#10000;
	data_in <= 24'b000011100001000000011000;
#10000;
	data_in <= 24'b000011000000111100010111;
#10000;
	data_in <= 24'b000010110000111000010110;
#10000;
	data_in <= 24'b000101010001100100101100;
#10000;
	data_in <= 24'b000101000001100000101010;
#10000;
	data_in <= 24'b000101010001100100101100;
#10000;
	data_in <= 24'b000101110001101100101101;
#10000;
	data_in <= 24'b000110000001110000101110;
#10000;
	data_in <= 24'b000101010001101000101001;
#10000;
	data_in <= 24'b000101010001101000101001;
#10000;
	data_in <= 24'b000101100001110000101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011001000100011000101101;
#10000;
	data_in <= 24'b010111100100001000101010;
#10000;
	data_in <= 24'b010111010100001000101101;
#10000;
	data_in <= 24'b011000010100100000110100;
#10000;
	data_in <= 24'b011000100100101000111000;
#10000;
	data_in <= 24'b010110110100010100110011;
#10000;
	data_in <= 24'b010011000011010100100101;
#10000;
	data_in <= 24'b001111000010010100010101;
#10000;
	data_in <= 24'b010100000011100100101001;
#10000;
	data_in <= 24'b010100100011111100110000;
#10000;
	data_in <= 24'b010111000100101100111110;
#10000;
	data_in <= 24'b010110100100101000111110;
#10000;
	data_in <= 24'b001111000010110100100100;
#10000;
	data_in <= 24'b000110100000110100000101;
#10000;
	data_in <= 24'b000011000000000000000000;
#10000;
	data_in <= 24'b000011100000001000000000;
#10000;
	data_in <= 24'b000100100000010100000011;
#10000;
	data_in <= 24'b000100100000100000001000;
#10000;
	data_in <= 24'b000101010000110100001110;
#10000;
	data_in <= 24'b000100110000111000010000;
#10000;
	data_in <= 24'b000010110000011100001100;
#10000;
	data_in <= 24'b000001010000010000001000;
#10000;
	data_in <= 24'b000001010000010100001011;
#10000;
	data_in <= 24'b000001110000011100001101;
#10000;
	data_in <= 24'b000011010000100000001010;
#10000;
	data_in <= 24'b000010010000100000001100;
#10000;
	data_in <= 24'b000010000000011000001100;
#10000;
	data_in <= 24'b000001000000001100001100;
#10000;
	data_in <= 24'b000000000000001000001010;
#10000;
	data_in <= 24'b000001000000011000010000;
#10000;
	data_in <= 24'b000000110000011100010010;
#10000;
	data_in <= 24'b000000000000001100001110;
#10000;
	data_in <= 24'b000010010000101100001011;
#10000;
	data_in <= 24'b000000110000010100000110;
#10000;
	data_in <= 24'b000001000000011000000111;
#10000;
	data_in <= 24'b000010100000101100001111;
#10000;
	data_in <= 24'b000001110000100000001100;
#10000;
	data_in <= 24'b000000010000010000001000;
#10000;
	data_in <= 24'b000000010000010000001001;
#10000;
	data_in <= 24'b000000110000011000001011;
#10000;
	data_in <= 24'b000011000001000000010001;
#10000;
	data_in <= 24'b000001100000101000001011;
#10000;
	data_in <= 24'b000001010000100000001100;
#10000;
	data_in <= 24'b000001110000101000001110;
#10000;
	data_in <= 24'b000001110000101000001110;
#10000;
	data_in <= 24'b000010010000110000010000;
#10000;
	data_in <= 24'b000010110000111000010010;
#10000;
	data_in <= 24'b000010100000110100010001;
#10000;
	data_in <= 24'b000010010000110000010100;
#10000;
	data_in <= 24'b000011010001001100011010;
#10000;
	data_in <= 24'b000100000001011000011011;
#10000;
	data_in <= 24'b000010110001000100010110;
#10000;
	data_in <= 24'b000001100000110000010001;
#10000;
	data_in <= 24'b000010010000111100010100;
#10000;
	data_in <= 24'b000010010001001000010110;
#10000;
	data_in <= 24'b000001010000111000010010;
#10000;
	data_in <= 24'b000110000001111000101011;
#10000;
	data_in <= 24'b000100000001011000100011;
#10000;
	data_in <= 24'b000011010001001100011110;
#10000;
	data_in <= 24'b000011110001010100100000;
#10000;
	data_in <= 24'b000011110001011000011111;
#10000;
	data_in <= 24'b000011110001011000011111;
#10000;
	data_in <= 24'b000011100001010100011110;
#10000;
	data_in <= 24'b000011000001001100011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001010110011001101010000;
#10000;
	data_in <= 24'b001110110100010101011101;
#10000;
	data_in <= 24'b001000100010110000111110;
#10000;
	data_in <= 24'b001101110100000101010011;
#10000;
	data_in <= 24'b010100110101101001110101;
#10000;
	data_in <= 24'b010001110100110101101010;
#10000;
	data_in <= 24'b010011110101011101110100;
#10000;
	data_in <= 24'b010100110110000001111010;
#10000;
	data_in <= 24'b000001010000111000110000;
#10000;
	data_in <= 24'b000100110001110100111011;
#10000;
	data_in <= 24'b000000000000110000100100;
#10000;
	data_in <= 24'b000000010000110100100101;
#10000;
	data_in <= 24'b000110010010000100111111;
#10000;
	data_in <= 24'b000111010010011001001000;
#10000;
	data_in <= 24'b001000100010101101010000;
#10000;
	data_in <= 24'b001000000011000001010101;
#10000;
	data_in <= 24'b000011100001010000110001;
#10000;
	data_in <= 24'b000101010001110100111010;
#10000;
	data_in <= 24'b000100000001101100110110;
#10000;
	data_in <= 24'b000010010001010000101111;
#10000;
	data_in <= 24'b000110010010001000111101;
#10000;
	data_in <= 24'b001001110010111101001101;
#10000;
	data_in <= 24'b001001000010101001001101;
#10000;
	data_in <= 24'b001000100010110001001110;
#10000;
	data_in <= 24'b000010110000110000100001;
#10000;
	data_in <= 24'b000010000000110100100010;
#10000;
	data_in <= 24'b000010110001001100101010;
#10000;
	data_in <= 24'b000010010001010000101010;
#10000;
	data_in <= 24'b000100000001100000101111;
#10000;
	data_in <= 24'b000101100001111000110101;
#10000;
	data_in <= 24'b000100010001010000110011;
#10000;
	data_in <= 24'b000100010001011000110101;
#10000;
	data_in <= 24'b000011100000100100010010;
#10000;
	data_in <= 24'b000001100000010100001111;
#10000;
	data_in <= 24'b000000000000010000010011;
#10000;
	data_in <= 24'b000000000000100100010111;
#10000;
	data_in <= 24'b000000000000011100010110;
#10000;
	data_in <= 24'b000000000000011000010101;
#10000;
	data_in <= 24'b000000100000010000011100;
#10000;
	data_in <= 24'b000000100000011000011110;
#10000;
	data_in <= 24'b000011110000100100001110;
#10000;
	data_in <= 24'b000011000000101000010000;
#10000;
	data_in <= 24'b000000100000011000010001;
#10000;
	data_in <= 24'b000000100000101000010111;
#10000;
	data_in <= 24'b000000100000100000010101;
#10000;
	data_in <= 24'b000001000000011100010110;
#10000;
	data_in <= 24'b000010110000110000100000;
#10000;
	data_in <= 24'b000001010000100000011101;
#10000;
	data_in <= 24'b000010110000010100010000;
#10000;
	data_in <= 24'b000010000000011000010010;
#10000;
	data_in <= 24'b000000100000100000010101;
#10000;
	data_in <= 24'b000001000000101100011010;
#10000;
	data_in <= 24'b000001110000101100011101;
#10000;
	data_in <= 24'b000010010000101000011110;
#10000;
	data_in <= 24'b000011100000110100100001;
#10000;
	data_in <= 24'b000010100000101100100000;
#10000;
	data_in <= 24'b000011100000100100011000;
#10000;
	data_in <= 24'b000001000000010000010010;
#10000;
	data_in <= 24'b000000000000010100010100;
#10000;
	data_in <= 24'b000000010000100000011001;
#10000;
	data_in <= 24'b000001100000011100011100;
#10000;
	data_in <= 24'b000001010000011000011011;
#10000;
	data_in <= 24'b000001100000010100011001;
#10000;
	data_in <= 24'b000010100000101100100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001110100100101101100110;
#10000;
	data_in <= 24'b001100010100011101100011;
#10000;
	data_in <= 24'b010100010110100110000111;
#10000;
	data_in <= 24'b001100100100110101101111;
#10000;
	data_in <= 24'b001011100100100001110000;
#10000;
	data_in <= 24'b001011100100100001110000;
#10000;
	data_in <= 24'b001100000100110101110100;
#10000;
	data_in <= 24'b001011110101001101110111;
#10000;
	data_in <= 24'b000110110011001101010111;
#10000;
	data_in <= 24'b000000000001110101000100;
#10000;
	data_in <= 24'b000111100011100101101011;
#10000;
	data_in <= 24'b001010110100011101111101;
#10000;
	data_in <= 24'b001011110100111010000001;
#10000;
	data_in <= 24'b001011110100111010000001;
#10000;
	data_in <= 24'b010000010110001010010100;
#10000;
	data_in <= 24'b001111100110011010010111;
#10000;
	data_in <= 24'b001001110011100101010110;
#10000;
	data_in <= 24'b001010110011111101011110;
#10000;
	data_in <= 24'b001010000011101101100001;
#10000;
	data_in <= 24'b001000100011010001011101;
#10000;
	data_in <= 24'b001010010011101001100001;
#10000;
	data_in <= 24'b001011100100000101100110;
#10000;
	data_in <= 24'b001110110101001001111000;
#10000;
	data_in <= 24'b001100110100110101110010;
#10000;
	data_in <= 24'b000010010001011100101110;
#10000;
	data_in <= 24'b000101100010011000111101;
#10000;
	data_in <= 24'b000011010001100000110110;
#10000;
	data_in <= 24'b000011000001011100110111;
#10000;
	data_in <= 24'b000100100001110000111010;
#10000;
	data_in <= 24'b000011000001100000110100;
#10000;
	data_in <= 24'b000011010001110000111100;
#10000;
	data_in <= 24'b000011010001111100111110;
#10000;
	data_in <= 24'b000000000000100000011100;
#10000;
	data_in <= 24'b000000000000010000011000;
#10000;
	data_in <= 24'b000000000000010100011100;
#10000;
	data_in <= 24'b000001110000111000100111;
#10000;
	data_in <= 24'b000001010000101000100011;
#10000;
	data_in <= 24'b000000000000100000100000;
#10000;
	data_in <= 24'b000000000000101000100110;
#10000;
	data_in <= 24'b000000000000110000100110;
#10000;
	data_in <= 24'b000000110000101000011110;
#10000;
	data_in <= 24'b000010110001010000101000;
#10000;
	data_in <= 24'b000100100001100100101101;
#10000;
	data_in <= 24'b000011000001001100100111;
#10000;
	data_in <= 24'b000011010000111100100111;
#10000;
	data_in <= 24'b000100110001100000110001;
#10000;
	data_in <= 24'b000100010001111100110110;
#10000;
	data_in <= 24'b000100100010000000110111;
#10000;
	data_in <= 24'b000001010000100100100101;
#10000;
	data_in <= 24'b000100100001100100110100;
#10000;
	data_in <= 24'b000101010001100100110101;
#10000;
	data_in <= 24'b000011100001001000101011;
#10000;
	data_in <= 24'b000100110001001000101100;
#10000;
	data_in <= 24'b000010100000101100100101;
#10000;
	data_in <= 24'b000001010000110000100101;
#10000;
	data_in <= 24'b000010100001010100110000;
#10000;
	data_in <= 24'b000010100000111000101010;
#10000;
	data_in <= 24'b000001100000110000101001;
#10000;
	data_in <= 24'b000001110000101100100111;
#10000;
	data_in <= 24'b000001110000101000100110;
#10000;
	data_in <= 24'b000010010000011100100100;
#10000;
	data_in <= 24'b000010110000100100100110;
#10000;
	data_in <= 24'b000101110001101100110111;
#10000;
	data_in <= 24'b000011100001010000110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001011110101110001111101;
#10000;
	data_in <= 24'b001101100110100110001010;
#10000;
	data_in <= 24'b001111000110110110010011;
#10000;
	data_in <= 24'b010010100111111010100110;
#10000;
	data_in <= 24'b010101011000101110110100;
#10000;
	data_in <= 24'b010111101001100111000001;
#10000;
	data_in <= 24'b010111001001101011000011;
#10000;
	data_in <= 24'b011000011010000111001010;
#10000;
	data_in <= 24'b001110100110101110011001;
#10000;
	data_in <= 24'b010000100111100010100111;
#10000;
	data_in <= 24'b010010000111110110110110;
#10000;
	data_in <= 24'b010011111000010111000001;
#10000;
	data_in <= 24'b010101101001001011001000;
#10000;
	data_in <= 24'b010111111010000011010011;
#10000;
	data_in <= 24'b011010111010110111100000;
#10000;
	data_in <= 24'b011110011011111011110000;
#10000;
	data_in <= 24'b010000100101111010000001;
#10000;
	data_in <= 24'b010001000110000010001001;
#10000;
	data_in <= 24'b010001010101111110010101;
#10000;
	data_in <= 24'b010000010101110010010101;
#10000;
	data_in <= 24'b010000100110000110010110;
#10000;
	data_in <= 24'b010000000110001010010111;
#10000;
	data_in <= 24'b010000110110101010011110;
#10000;
	data_in <= 24'b010010000111001010100111;
#10000;
	data_in <= 24'b000000010001000100101110;
#10000;
	data_in <= 24'b000000110000111100110001;
#10000;
	data_in <= 24'b000001010000111100111110;
#10000;
	data_in <= 24'b000000000000101100111101;
#10000;
	data_in <= 24'b000001000001010001000011;
#10000;
	data_in <= 24'b000000000001001001000001;
#10000;
	data_in <= 24'b000000010001011101000111;
#10000;
	data_in <= 24'b000000000001100101001000;
#10000;
	data_in <= 24'b000001100001001000101010;
#10000;
	data_in <= 24'b000001110001000000101011;
#10000;
	data_in <= 24'b000010100001001100110100;
#10000;
	data_in <= 24'b000001100000111100110100;
#10000;
	data_in <= 24'b000010000001011000111010;
#10000;
	data_in <= 24'b000001100001100000111101;
#10000;
	data_in <= 24'b000100000010001101001000;
#10000;
	data_in <= 24'b000100100010011101001101;
#10000;
	data_in <= 24'b000110000010000000110111;
#10000;
	data_in <= 24'b000101100001110000110011;
#10000;
	data_in <= 24'b000101000001101100110110;
#10000;
	data_in <= 24'b000011100001100100110101;
#10000;
	data_in <= 24'b000011000001011100110111;
#10000;
	data_in <= 24'b000010110001011100111001;
#10000;
	data_in <= 24'b000011100001110100111110;
#10000;
	data_in <= 24'b000011010001110000111101;
#10000;
	data_in <= 24'b000010100001000000101101;
#10000;
	data_in <= 24'b000010010000111100101100;
#10000;
	data_in <= 24'b000011000001001100101100;
#10000;
	data_in <= 24'b000011100001011100110010;
#10000;
	data_in <= 24'b000010110001001000110011;
#10000;
	data_in <= 24'b000011100001010000110111;
#10000;
	data_in <= 24'b000011010001001100110110;
#10000;
	data_in <= 24'b000010100001000000110011;
#10000;
	data_in <= 24'b000001000000100100101010;
#10000;
	data_in <= 24'b000010110001000000101111;
#10000;
	data_in <= 24'b000100100001100100110100;
#10000;
	data_in <= 24'b000101100001110100111000;
#10000;
	data_in <= 24'b000001110000110000101101;
#10000;
	data_in <= 24'b000010010000110100110000;
#10000;
	data_in <= 24'b000011000001000000110011;
#10000;
	data_in <= 24'b000100000001010000110111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b011000011010001011001001;
#10000;
	data_in <= 24'b011010001010100111010000;
#10000;
	data_in <= 24'b011010111010101011010000;
#10000;
	data_in <= 24'b011100111010111111010011;
#10000;
	data_in <= 24'b100000001011011111011100;
#10000;
	data_in <= 24'b100010011011111011011111;
#10000;
	data_in <= 24'b100101101100100011100110;
#10000;
	data_in <= 24'b100111001100111011100101;
#10000;
	data_in <= 24'b011111001100000111110010;
#10000;
	data_in <= 24'b100010101101000111111101;
#10000;
	data_in <= 24'b100100111101100011111111;
#10000;
	data_in <= 24'b100111011101111011111111;
#10000;
	data_in <= 24'b101010001110010011111111;
#10000;
	data_in <= 24'b101011101110101011111111;
#10000;
	data_in <= 24'b101101111111000111111111;
#10000;
	data_in <= 24'b101110011111000111111111;
#10000;
	data_in <= 24'b010001100111010110101000;
#10000;
	data_in <= 24'b010100101000001110110101;
#10000;
	data_in <= 24'b010101101000101110111101;
#10000;
	data_in <= 24'b010111111001011011001001;
#10000;
	data_in <= 24'b011001111001110111011001;
#10000;
	data_in <= 24'b011010101010001111011011;
#10000;
	data_in <= 24'b011100011010110111011011;
#10000;
	data_in <= 24'b011100111011000111011010;
#10000;
	data_in <= 24'b000001100010010001010011;
#10000;
	data_in <= 24'b000001100010101001011010;
#10000;
	data_in <= 24'b000001010010110101011101;
#10000;
	data_in <= 24'b000011110011101001101101;
#10000;
	data_in <= 24'b000101000100000001111101;
#10000;
	data_in <= 24'b000100100100000101111110;
#10000;
	data_in <= 24'b000110000100110110000000;
#10000;
	data_in <= 24'b001000000101010110000111;
#10000;
	data_in <= 24'b000011100010100001001101;
#10000;
	data_in <= 24'b000100000010101101010000;
#10000;
	data_in <= 24'b000011000010100101010000;
#10000;
	data_in <= 24'b000100000010110101011001;
#10000;
	data_in <= 24'b000101010011000001100010;
#10000;
	data_in <= 24'b000100110011000001100011;
#10000;
	data_in <= 24'b000101010011010001100111;
#10000;
	data_in <= 24'b000110100011011101101010;
#10000;
	data_in <= 24'b000010110001110000111101;
#10000;
	data_in <= 24'b000100000010001101000100;
#10000;
	data_in <= 24'b000010110001111001000001;
#10000;
	data_in <= 24'b000010000001101000111111;
#10000;
	data_in <= 24'b000010100001110101000011;
#10000;
	data_in <= 24'b000011110010001001001101;
#10000;
	data_in <= 24'b000101010010011001010111;
#10000;
	data_in <= 24'b000100110010010001010111;
#10000;
	data_in <= 24'b000011100001010100110110;
#10000;
	data_in <= 24'b000100110001110000111101;
#10000;
	data_in <= 24'b000100010001101000111011;
#10000;
	data_in <= 24'b000011110001101000111010;
#10000;
	data_in <= 24'b000011100001110100111101;
#10000;
	data_in <= 24'b000011110001111101000011;
#10000;
	data_in <= 24'b000101000010001101010001;
#10000;
	data_in <= 24'b000101000010010101011000;
#10000;
	data_in <= 24'b000100010001011000110111;
#10000;
	data_in <= 24'b000101010001101000111011;
#10000;
	data_in <= 24'b000101110001111000111111;
#10000;
	data_in <= 24'b000111110010100001001001;
#10000;
	data_in <= 24'b000111000010011101000111;
#10000;
	data_in <= 24'b000010110001100100111101;
#10000;
	data_in <= 24'b000010110001100001000110;
#10000;
	data_in <= 24'b000100010001111101010000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b101010011101110111101110;
#10000;
	data_in <= 24'b101111101110101011111011;
#10000;
	data_in <= 24'b110011011110100111111111;
#10000;
	data_in <= 24'b010000110101000001101010;
#10000;
	data_in <= 24'b000101000001010000101100;
#10000;
	data_in <= 24'b011111000111101010001110;
#10000;
	data_in <= 24'b110010111100111111100001;
#10000;
	data_in <= 24'b110110101110100111111001;
#10000;
	data_in <= 24'b110000001111011011111111;
#10000;
	data_in <= 24'b110001101111011111111111;
#10000;
	data_in <= 24'b110100001111011111111111;
#10000;
	data_in <= 24'b100100111011000011001111;
#10000;
	data_in <= 24'b001100100100011001100101;
#10000;
	data_in <= 24'b100110001010101111000110;
#10000;
	data_in <= 24'b110111101111010111111111;
#10000;
	data_in <= 24'b110110101111101011111111;
#10000;
	data_in <= 24'b011110011011001011011111;
#10000;
	data_in <= 24'b011111001011001011100001;
#10000;
	data_in <= 24'b011111011011000111100000;
#10000;
	data_in <= 24'b100111101100111111111111;
#10000;
	data_in <= 24'b100001101011001011100001;
#10000;
	data_in <= 24'b100101011100001011101101;
#10000;
	data_in <= 24'b100110001100100011110010;
#10000;
	data_in <= 24'b101000011101100011111111;
#10000;
	data_in <= 24'b000111110100111010000110;
#10000;
	data_in <= 24'b001110000110011110011111;
#10000;
	data_in <= 24'b001100110110010110011111;
#10000;
	data_in <= 24'b001100110110011010011110;
#10000;
	data_in <= 24'b001101010110011110011100;
#10000;
	data_in <= 24'b001100110110010110011010;
#10000;
	data_in <= 24'b010000110111101010101101;
#10000;
	data_in <= 24'b010001111000010010110110;
#10000;
	data_in <= 24'b000110010011010101101011;
#10000;
	data_in <= 24'b000110010011010101101011;
#10000;
	data_in <= 24'b000101110011011001101101;
#10000;
	data_in <= 24'b000111110100001101111001;
#10000;
	data_in <= 24'b001010000100101010000000;
#10000;
	data_in <= 24'b001001100100101110000011;
#10000;
	data_in <= 24'b001110000110000010011010;
#10000;
	data_in <= 24'b001110110110101110100101;
#10000;
	data_in <= 24'b000100000010001101010110;
#10000;
	data_in <= 24'b000110110011000001100011;
#10000;
	data_in <= 24'b001000010011100001101010;
#10000;
	data_in <= 24'b000111010011010101101001;
#10000;
	data_in <= 24'b001001100011111001110100;
#10000;
	data_in <= 24'b001001010011111001110110;
#10000;
	data_in <= 24'b001011000100100010000100;
#10000;
	data_in <= 24'b001100110101011110010011;
#10000;
	data_in <= 24'b000100010010010001010111;
#10000;
	data_in <= 24'b000100010010011101010111;
#10000;
	data_in <= 24'b000111000011001101100011;
#10000;
	data_in <= 24'b000110010010111101011111;
#10000;
	data_in <= 24'b000111110011000001100011;
#10000;
	data_in <= 24'b000111110010111101100100;
#10000;
	data_in <= 24'b001010000011101101110100;
#10000;
	data_in <= 24'b001000010011110001110100;
#10000;
	data_in <= 24'b000101000010010101010110;
#10000;
	data_in <= 24'b000101100010101001011010;
#10000;
	data_in <= 24'b000001100001101001001010;
#10000;
	data_in <= 24'b000011000001110101001110;
#10000;
	data_in <= 24'b000011010001101101001111;
#10000;
	data_in <= 24'b000100100010000001010101;
#10000;
	data_in <= 24'b000010000001100101010001;
#10000;
	data_in <= 24'b000010010010000001011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b110101101111001011111111;
#10000;
	data_in <= 24'b110001111110100111111001;
#10000;
	data_in <= 24'b110101001111010111111111;
#10000;
	data_in <= 24'b110111111111110011111111;
#10000;
	data_in <= 24'b111000111111110111111111;
#10000;
	data_in <= 24'b110111111111100111111111;
#10000;
	data_in <= 24'b110010011110101011111101;
#10000;
	data_in <= 24'b110000111110110011111111;
#10000;
	data_in <= 24'b110011111111101111111111;
#10000;
	data_in <= 24'b101001001101011011101100;
#10000;
	data_in <= 24'b101011111110000011110110;
#10000;
	data_in <= 24'b101100111110001011110111;
#10000;
	data_in <= 24'b101101111110001011110111;
#10000;
	data_in <= 24'b101001011100111111100110;
#10000;
	data_in <= 24'b100001001011001111001111;
#10000;
	data_in <= 24'b010110101001000010101111;
#10000;
	data_in <= 24'b100110101101101111111111;
#10000;
	data_in <= 24'b100001001100101011101111;
#10000;
	data_in <= 24'b100011011101001111111000;
#10000;
	data_in <= 24'b100011001101000011110011;
#10000;
	data_in <= 24'b100110101101101011111101;
#10000;
	data_in <= 24'b100100001101000011110011;
#10000;
	data_in <= 24'b011111001100001011100111;
#10000;
	data_in <= 24'b011011011011011011011100;
#10000;
	data_in <= 24'b010010111001000011000010;
#10000;
	data_in <= 24'b010111001010100011011001;
#10000;
	data_in <= 24'b011101111100010011110101;
#10000;
	data_in <= 24'b100001101101001011111111;
#10000;
	data_in <= 24'b100011111101100111111111;
#10000;
	data_in <= 24'b100011011101011111111111;
#10000;
	data_in <= 24'b011111101100110011111011;
#10000;
	data_in <= 24'b011111011100110111111100;
#10000;
	data_in <= 24'b010001000111110110111010;
#10000;
	data_in <= 24'b010001111000100011000101;
#10000;
	data_in <= 24'b010110101001110111011100;
#10000;
	data_in <= 24'b011000011010011011100101;
#10000;
	data_in <= 24'b010111101010000111100000;
#10000;
	data_in <= 24'b011000011010011111100011;
#10000;
	data_in <= 24'b010100111010000011011001;
#10000;
	data_in <= 24'b010000111000110011000110;
#10000;
	data_in <= 24'b001011100101110110011011;
#10000;
	data_in <= 24'b001101010110101110101010;
#10000;
	data_in <= 24'b010010111000001111000100;
#10000;
	data_in <= 24'b010011011000011111001001;
#10000;
	data_in <= 24'b010110101001001111011000;
#10000;
	data_in <= 24'b010100111000111011010011;
#10000;
	data_in <= 24'b010001101000100011001001;
#10000;
	data_in <= 24'b001101010111001110110011;
#10000;
	data_in <= 24'b000100110011101101110000;
#10000;
	data_in <= 24'b001001000101001010001000;
#10000;
	data_in <= 24'b001101100110001010011101;
#10000;
	data_in <= 24'b001101100110000110100000;
#10000;
	data_in <= 24'b010010000110111110110011;
#10000;
	data_in <= 24'b001101010101111010100011;
#10000;
	data_in <= 24'b001001010101011010011010;
#10000;
	data_in <= 24'b001000010101001110010101;
#10000;
	data_in <= 24'b000001100010011001011011;
#10000;
	data_in <= 24'b000010110010111101100101;
#10000;
	data_in <= 24'b000110110011110101111000;
#10000;
	data_in <= 24'b001100000100111110001100;
#10000;
	data_in <= 24'b001101000101001010010011;
#10000;
	data_in <= 24'b001011100100111010010000;
#10000;
	data_in <= 24'b001001000100100110001101;
#10000;
	data_in <= 24'b000111100100010010000101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b100111001100110011101000;
#10000;
	data_in <= 24'b100010111011111111011101;
#10000;
	data_in <= 24'b100011111100000111011111;
#10000;
	data_in <= 24'b011101101010101011001000;
#10000;
	data_in <= 24'b011111011011011111010100;
#10000;
	data_in <= 24'b100010101100101011101000;
#10000;
	data_in <= 24'b011001011010100011000111;
#10000;
	data_in <= 24'b010111101001110110111111;
#10000;
	data_in <= 24'b011000111010001111000010;
#10000;
	data_in <= 24'b011111111100010011100101;
#10000;
	data_in <= 24'b101001001110101111111111;
#10000;
	data_in <= 24'b101000011110101011111111;
#10000;
	data_in <= 24'b100100111110001011111111;
#10000;
	data_in <= 24'b100011001101111011111111;
#10000;
	data_in <= 24'b011101101100011111101100;
#10000;
	data_in <= 24'b011100101011110011100110;
#10000;
	data_in <= 24'b011101001100000111101000;
#10000;
	data_in <= 24'b100000111101001111111100;
#10000;
	data_in <= 24'b100011101110000111111111;
#10000;
	data_in <= 24'b100011101110001111111111;
#10000;
	data_in <= 24'b100000011101110011111111;
#10000;
	data_in <= 24'b011110111101010111111110;
#10000;
	data_in <= 24'b011111011101001011111111;
#10000;
	data_in <= 24'b011110111100100011111001;
#10000;
	data_in <= 24'b011010101011011011100111;
#10000;
	data_in <= 24'b011000011010110111011101;
#10000;
	data_in <= 24'b010101111010001111010011;
#10000;
	data_in <= 24'b010101101010010011010010;
#10000;
	data_in <= 24'b010010011001101011000111;
#10000;
	data_in <= 24'b001111011000110110111100;
#10000;
	data_in <= 24'b010000011000110110111110;
#10000;
	data_in <= 24'b010000101000011010111011;
#10000;
	data_in <= 24'b001101010111000110101100;
#10000;
	data_in <= 24'b001010110101111110011011;
#10000;
	data_in <= 24'b001001010101100010010000;
#10000;
	data_in <= 24'b001001110101100110001110;
#10000;
	data_in <= 24'b001000110101100010001011;
#10000;
	data_in <= 24'b000111110101010010000111;
#10000;
	data_in <= 24'b000111110100111110000011;
#10000;
	data_in <= 24'b000110110100011101111100;
#10000;
	data_in <= 24'b001101010110010110100101;
#10000;
	data_in <= 24'b001011000101001010010010;
#10000;
	data_in <= 24'b001001010100011010000101;
#10000;
	data_in <= 24'b000111110011110101111000;
#10000;
	data_in <= 24'b001000000011111101110110;
#10000;
	data_in <= 24'b001001000100010001111001;
#10000;
	data_in <= 24'b000110010011100001101011;
#10000;
	data_in <= 24'b000100000010111001011111;
#10000;
	data_in <= 24'b000011000011011001110111;
#10000;
	data_in <= 24'b000100110011010001110011;
#10000;
	data_in <= 24'b000111000011001101110001;
#10000;
	data_in <= 24'b000111100011000001101011;
#10000;
	data_in <= 24'b000110110010111101100110;
#10000;
	data_in <= 24'b000101010010101001011101;
#10000;
	data_in <= 24'b000011000010010001010010;
#10000;
	data_in <= 24'b000011000010001101010000;
#10000;
	data_in <= 24'b000110100011110101111101;
#10000;
	data_in <= 24'b000101110011001101110000;
#10000;
	data_in <= 24'b000100010010010001100001;
#10000;
	data_in <= 24'b000101110010010101011111;
#10000;
	data_in <= 24'b000101100010010001011001;
#10000;
	data_in <= 24'b000010010001100001001001;
#10000;
	data_in <= 24'b000010000001101001001001;
#10000;
	data_in <= 24'b000101000010011101010010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001101100110101010001111;
#10000;
	data_in <= 24'b000000000001100101000000;
#10000;
	data_in <= 24'b000000110010011001001110;
#10000;
	data_in <= 24'b000000000001111101000110;
#10000;
	data_in <= 24'b000000000001010100111000;
#10000;
	data_in <= 24'b000000000001000000110001;
#10000;
	data_in <= 24'b000000000000111000101101;
#10000;
	data_in <= 24'b000001110010001101000010;
#10000;
	data_in <= 24'b011011111010101111011001;
#10000;
	data_in <= 24'b010110011000111011000000;
#10000;
	data_in <= 24'b010111111000111111000011;
#10000;
	data_in <= 24'b010111111000111011000001;
#10000;
	data_in <= 24'b011001001001001111000110;
#10000;
	data_in <= 24'b011000101001000011000000;
#10000;
	data_in <= 24'b011010011000111110111111;
#10000;
	data_in <= 24'b010110110111111110101111;
#10000;
	data_in <= 24'b011110111011110011110011;
#10000;
	data_in <= 24'b011101101011000011101011;
#10000;
	data_in <= 24'b011000011001101011010111;
#10000;
	data_in <= 24'b010101011000111011001011;
#10000;
	data_in <= 24'b010110001001000111001110;
#10000;
	data_in <= 24'b010011001000001010111110;
#10000;
	data_in <= 24'b010101011000000110111110;
#10000;
	data_in <= 24'b010001010110110110100111;
#10000;
	data_in <= 24'b001111010111010110110000;
#10000;
	data_in <= 24'b001110010110110010101010;
#10000;
	data_in <= 24'b001101100110100110100111;
#10000;
	data_in <= 24'b001011000110000110100000;
#10000;
	data_in <= 24'b001011110110010110100010;
#10000;
	data_in <= 24'b001011110110000010011110;
#10000;
	data_in <= 24'b001110000101111010011110;
#10000;
	data_in <= 24'b001110100101111010011010;
#10000;
	data_in <= 24'b001000000100001101111011;
#10000;
	data_in <= 24'b000111100011111101110111;
#10000;
	data_in <= 24'b001001100100011101111111;
#10000;
	data_in <= 24'b000101000011010101101101;
#10000;
	data_in <= 24'b000010100010111001100100;
#10000;
	data_in <= 24'b000100110011001101101000;
#10000;
	data_in <= 24'b000101110010111101100101;
#10000;
	data_in <= 24'b000100010010011101011011;
#10000;
	data_in <= 24'b000100010010100001011010;
#10000;
	data_in <= 24'b000011110010010001010111;
#10000;
	data_in <= 24'b000100010010011001011001;
#10000;
	data_in <= 24'b000011000010001101010011;
#10000;
	data_in <= 24'b000001110001111001001110;
#10000;
	data_in <= 24'b000100000010011101010101;
#10000;
	data_in <= 24'b000111110010111001011100;
#10000;
	data_in <= 24'b000100010010000101001100;
#10000;
	data_in <= 24'b000100010010010001010001;
#10000;
	data_in <= 24'b000011100001111001001100;
#10000;
	data_in <= 24'b000011010001111001001001;
#10000;
	data_in <= 24'b000101010010011101010000;
#10000;
	data_in <= 24'b000100010010010101001110;
#10000;
	data_in <= 24'b000011110010001001001000;
#10000;
	data_in <= 24'b000101000010010001001001;
#10000;
	data_in <= 24'b000011100001101000111110;
#10000;
	data_in <= 24'b000101000010010001001111;
#10000;
	data_in <= 24'b000100100010000001001010;
#10000;
	data_in <= 24'b000100110010000101001011;
#10000;
	data_in <= 24'b000100110010001001001001;
#10000;
	data_in <= 24'b000100100010001001000111;
#10000;
	data_in <= 24'b000101000010010001001000;
#10000;
	data_in <= 24'b000011110001111000111111;
#10000;
	data_in <= 24'b000101000001111001000000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000010010010001101000111;
#10000;
	data_in <= 24'b000100100010100101001111;
#10000;
	data_in <= 24'b000100010010100001001110;
#10000;
	data_in <= 24'b001000010011100001011110;
#10000;
	data_in <= 24'b000110000010111001010010;
#10000;
	data_in <= 24'b001000000011011001011010;
#10000;
	data_in <= 24'b001010110100000101100101;
#10000;
	data_in <= 24'b001100110100100101101101;
#10000;
	data_in <= 24'b010010110110111110011111;
#10000;
	data_in <= 24'b010010110110111010100000;
#10000;
	data_in <= 24'b010000000110001110010101;
#10000;
	data_in <= 24'b010000100110001110010100;
#10000;
	data_in <= 24'b010000000110000110010010;
#10000;
	data_in <= 24'b001110000101101010001000;
#10000;
	data_in <= 24'b001110100101101110001001;
#10000;
	data_in <= 24'b001111100101110010001011;
#10000;
	data_in <= 24'b010001110111000110100110;
#10000;
	data_in <= 24'b010001010110110110100001;
#10000;
	data_in <= 24'b001101110101111110010011;
#10000;
	data_in <= 24'b001011010101010110000110;
#10000;
	data_in <= 24'b001110110110000010010010;
#10000;
	data_in <= 24'b001011010101000110000001;
#10000;
	data_in <= 24'b001010100100110001111010;
#10000;
	data_in <= 24'b001010010100101001110111;
#10000;
	data_in <= 24'b001101110101110110010011;
#10000;
	data_in <= 24'b001100000101100010001001;
#10000;
	data_in <= 24'b001001100100111001111111;
#10000;
	data_in <= 24'b000111000100001001110010;
#10000;
	data_in <= 24'b001001110100101101111011;
#10000;
	data_in <= 24'b000110110011110101101011;
#10000;
	data_in <= 24'b000101100011100001100011;
#10000;
	data_in <= 24'b000101110011010101011110;
#10000;
	data_in <= 24'b000101000011000001011111;
#10000;
	data_in <= 24'b000011010010110001011001;
#10000;
	data_in <= 24'b000011110010111001011011;
#10000;
	data_in <= 24'b000100000010110101011001;
#10000;
	data_in <= 24'b000011110010110001011000;
#10000;
	data_in <= 24'b000100010010110101010110;
#10000;
	data_in <= 24'b000101000010111001010110;
#10000;
	data_in <= 24'b000101100010110101010011;
#10000;
	data_in <= 24'b000011100001111101001010;
#10000;
	data_in <= 24'b000010100001111001000111;
#10000;
	data_in <= 24'b000011100010001001001011;
#10000;
	data_in <= 24'b000100100010010101001011;
#10000;
	data_in <= 24'b000010000001101101000001;
#10000;
	data_in <= 24'b000011000001111101000101;
#10000;
	data_in <= 24'b000011000001111001000011;
#10000;
	data_in <= 24'b000011010010000001000011;
#10000;
	data_in <= 24'b000100010001100100111110;
#10000;
	data_in <= 24'b000101000001101000111111;
#10000;
	data_in <= 24'b000110000001111001000011;
#10000;
	data_in <= 24'b000101110001111101000100;
#10000;
	data_in <= 24'b000101100001111001000011;
#10000;
	data_in <= 24'b000110100010001101001000;
#10000;
	data_in <= 24'b000101000001110101000010;
#10000;
	data_in <= 24'b000110000010001001000100;
#10000;
	data_in <= 24'b000101100001101100111100;
#10000;
	data_in <= 24'b000110100001101100111101;
#10000;
	data_in <= 24'b000101110001100100111011;
#10000;
	data_in <= 24'b000100100001010000110110;
#10000;
	data_in <= 24'b000110000001110100111110;
#10000;
	data_in <= 24'b000101110001110000111101;
#10000;
	data_in <= 24'b000001100000110100101110;
#10000;
	data_in <= 24'b000010110001001000110011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b001000000011001101011000;
#10000;
	data_in <= 24'b000101110010101001001111;
#10000;
	data_in <= 24'b000001110001101000111111;
#10000;
	data_in <= 24'b000110000010101101010000;
#10000;
	data_in <= 24'b000110110010111001010011;
#10000;
	data_in <= 24'b001001100011100101011110;
#10000;
	data_in <= 24'b000111110011001001010111;
#10000;
	data_in <= 24'b000111000010111101010010;
#10000;
	data_in <= 24'b001111000101100110000110;
#10000;
	data_in <= 24'b001100100100110001111010;
#10000;
	data_in <= 24'b001001110011111101101101;
#10000;
	data_in <= 24'b001010010100001001101110;
#10000;
	data_in <= 24'b001001010011111001101010;
#10000;
	data_in <= 24'b001010010100000001101101;
#10000;
	data_in <= 24'b001010010100000001101101;
#10000;
	data_in <= 24'b001000010011011101100000;
#10000;
	data_in <= 24'b001011100100101101110111;
#10000;
	data_in <= 24'b001011100100011101110001;
#10000;
	data_in <= 24'b001010100100001101101011;
#10000;
	data_in <= 24'b001000100011100101011111;
#10000;
	data_in <= 24'b000111000011001001010110;
#10000;
	data_in <= 24'b000100110010011001001011;
#10000;
	data_in <= 24'b000100000010001101000110;
#10000;
	data_in <= 24'b000000110001010000110101;
#10000;
	data_in <= 24'b000101100011000001011000;
#10000;
	data_in <= 24'b001001010011110001100010;
#10000;
	data_in <= 24'b000100010010010101001000;
#10000;
	data_in <= 24'b000000000001000000110001;
#10000;
	data_in <= 24'b000010100001110000111011;
#10000;
	data_in <= 24'b000010000001100000110101;
#10000;
	data_in <= 24'b000001110001010100110001;
#10000;
	data_in <= 24'b000101100010001000111110;
#10000;
	data_in <= 24'b000011110010010101001000;
#10000;
	data_in <= 24'b000100010010010001000101;
#10000;
	data_in <= 24'b000110010010100101000110;
#10000;
	data_in <= 24'b000111110010110101001001;
#10000;
	data_in <= 24'b000101100010001000111010;
#10000;
	data_in <= 24'b000111000010011100111101;
#10000;
	data_in <= 24'b001000100010110101000011;
#10000;
	data_in <= 24'b000101000001111000110110;
#10000;
	data_in <= 24'b000100110010001001000011;
#10000;
	data_in <= 24'b000111100010110001001001;
#10000;
	data_in <= 24'b000110000010010001000000;
#10000;
	data_in <= 24'b000110100010010101000000;
#10000;
	data_in <= 24'b000111100010100001000000;
#10000;
	data_in <= 24'b000111010010010100111100;
#10000;
	data_in <= 24'b000110000010000100110101;
#10000;
	data_in <= 24'b000110100010001000111001;
#10000;
	data_in <= 24'b000100100001110100111101;
#10000;
	data_in <= 24'b000100010001110000111100;
#10000;
	data_in <= 24'b000011110001100100110111;
#10000;
	data_in <= 24'b000100010001110000111000;
#10000;
	data_in <= 24'b000110000010000100111100;
#10000;
	data_in <= 24'b000100010001101000110101;
#10000;
	data_in <= 24'b000101010001111100110111;
#10000;
	data_in <= 24'b000110000001111100111000;
#10000;
	data_in <= 24'b000011110001011100110101;
#10000;
	data_in <= 24'b000000010000101100101001;
#10000;
	data_in <= 24'b000010110001001100110000;
#10000;
	data_in <= 24'b000011100001011000110011;
#10000;
	data_in <= 24'b000100000001100000110101;
#10000;
	data_in <= 24'b000001010000110000100111;
#10000;
	data_in <= 24'b000100000001011100110010;
#10000;
	data_in <= 24'b000010100001000100101010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000110110010110101001010;
#10000;
	data_in <= 24'b000111110011000001001010;
#10000;
	data_in <= 24'b001000110011000101001101;
#10000;
	data_in <= 24'b000111000010101101000101;
#10000;
	data_in <= 24'b000111100010101101000101;
#10000;
	data_in <= 24'b000110010010011100111110;
#10000;
	data_in <= 24'b000101100010001000111010;
#10000;
	data_in <= 24'b000011110001101000110000;
#10000;
	data_in <= 24'b001000100011011101010111;
#10000;
	data_in <= 24'b001000100011011001010101;
#10000;
	data_in <= 24'b001000010011010101010100;
#10000;
	data_in <= 24'b000111100011000001001111;
#10000;
	data_in <= 24'b000111100011000001001101;
#10000;
	data_in <= 24'b001000000011000001001101;
#10000;
	data_in <= 24'b000110110010110001000111;
#10000;
	data_in <= 24'b000100100010000000111100;
#10000;
	data_in <= 24'b000001000001001100110011;
#10000;
	data_in <= 24'b000001100001010000110001;
#10000;
	data_in <= 24'b000010010001011100110100;
#10000;
	data_in <= 24'b000010100001100000110101;
#10000;
	data_in <= 24'b000010110001100100110110;
#10000;
	data_in <= 24'b000100110010001101000000;
#10000;
	data_in <= 24'b000101010010011001000001;
#10000;
	data_in <= 24'b000011000001110100111000;
#10000;
	data_in <= 24'b000011010001100000110110;
#10000;
	data_in <= 24'b000100000001101100111001;
#10000;
	data_in <= 24'b000100110001111000111100;
#10000;
	data_in <= 24'b000100010001110000111010;
#10000;
	data_in <= 24'b000010010001010000110010;
#10000;
	data_in <= 24'b000011010001101100111000;
#10000;
	data_in <= 24'b000100010001111100111011;
#10000;
	data_in <= 24'b000011000001101000110110;
#10000;
	data_in <= 24'b000101000001111100111011;
#10000;
	data_in <= 24'b000101100010000100111111;
#10000;
	data_in <= 24'b000110110010011001000100;
#10000;
	data_in <= 24'b000110110010011001000100;
#10000;
	data_in <= 24'b000110000010001101000001;
#10000;
	data_in <= 24'b000111010010011101000101;
#10000;
	data_in <= 24'b001000100010110001001010;
#10000;
	data_in <= 24'b001000000010101001001000;
#10000;
	data_in <= 24'b000110010010001000111101;
#10000;
	data_in <= 24'b000101000001111100111011;
#10000;
	data_in <= 24'b000101000001111100111011;
#10000;
	data_in <= 24'b000100000001101100110111;
#10000;
	data_in <= 24'b000101000001111100111011;
#10000;
	data_in <= 24'b000100000001100000110101;
#10000;
	data_in <= 24'b000100000001100000110101;
#10000;
	data_in <= 24'b000011010001010100110010;
#10000;
	data_in <= 24'b000101110001111100110110;
#10000;
	data_in <= 24'b000100110001100100110000;
#10000;
	data_in <= 24'b000100100001101000110001;
#10000;
	data_in <= 24'b000010100001001000101001;
#10000;
	data_in <= 24'b000110000010000000110111;
#10000;
	data_in <= 24'b000010010001010000101010;
#10000;
	data_in <= 24'b000010100001010000101100;
#10000;
	data_in <= 24'b000011000001011000101110;
#10000;
	data_in <= 24'b000011000001000100100110;
#10000;
	data_in <= 24'b000010100001000000100011;
#10000;
	data_in <= 24'b000011100001001100101000;
#10000;
	data_in <= 24'b000001100000110100100001;
#10000;
	data_in <= 24'b000110100010000100110101;
#10000;
	data_in <= 24'b000010100001000100100101;
#10000;
	data_in <= 24'b000011110001011100101110;
#10000;
	data_in <= 24'b000110000010000000110111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000101100001111000110101;
#10000;
	data_in <= 24'b000101000001101100101111;
#10000;
	data_in <= 24'b000110100010000100110100;
#10000;
	data_in <= 24'b000110100010000000110011;
#10000;
	data_in <= 24'b000011100001001000100100;
#10000;
	data_in <= 24'b000011100001001000100100;
#10000;
	data_in <= 24'b000110010001101100101101;
#10000;
	data_in <= 24'b000101110001100100101011;
#10000;
	data_in <= 24'b000110000010010100111111;
#10000;
	data_in <= 24'b000110110010011001000001;
#10000;
	data_in <= 24'b000011110001100100110001;
#10000;
	data_in <= 24'b000011000001010000101011;
#10000;
	data_in <= 24'b000110110010001000110110;
#10000;
	data_in <= 24'b000110010001111000110011;
#10000;
	data_in <= 24'b000011110001010000101001;
#10000;
	data_in <= 24'b000101010001100000101101;
#10000;
	data_in <= 24'b000100000001111100111001;
#10000;
	data_in <= 24'b000100100010000100111011;
#10000;
	data_in <= 24'b000010110001101100110010;
#10000;
	data_in <= 24'b000011000001101000110000;
#10000;
	data_in <= 24'b000101010010010000110111;
#10000;
	data_in <= 24'b000101000010001000110101;
#10000;
	data_in <= 24'b000011000001101000101101;
#10000;
	data_in <= 24'b000011010001101100101110;
#10000;
	data_in <= 24'b000100100010000000111100;
#10000;
	data_in <= 24'b000100000001111100111001;
#10000;
	data_in <= 24'b000100010001111000111000;
#10000;
	data_in <= 24'b000011100001110000110011;
#10000;
	data_in <= 24'b000010100001011100101101;
#10000;
	data_in <= 24'b000010000001010100101011;
#10000;
	data_in <= 24'b000001110001010000101010;
#10000;
	data_in <= 24'b000001100001010000100111;
#10000;
	data_in <= 24'b000110000010000000111110;
#10000;
	data_in <= 24'b000101110001111100111100;
#10000;
	data_in <= 24'b000100000001011000110011;
#10000;
	data_in <= 24'b000010100001000100101100;
#10000;
	data_in <= 24'b000011110001001100101111;
#10000;
	data_in <= 24'b000011100001001100101100;
#10000;
	data_in <= 24'b000011010001000100101010;
#10000;
	data_in <= 24'b000100010001010100101101;
#10000;
	data_in <= 24'b000100100001100000110101;
#10000;
	data_in <= 24'b000011100001010000110001;
#10000;
	data_in <= 24'b000100010001010100110001;
#10000;
	data_in <= 24'b000100110001011000110010;
#10000;
	data_in <= 24'b000100100001011000101111;
#10000;
	data_in <= 24'b000101000001100000110001;
#10000;
	data_in <= 24'b000110000001101000110010;
#10000;
	data_in <= 24'b000101100001100000110000;
#10000;
	data_in <= 24'b000010110001010100101101;
#10000;
	data_in <= 24'b000011000001001100101100;
#10000;
	data_in <= 24'b000101010001110100110100;
#10000;
	data_in <= 24'b000110010001111100110110;
#10000;
	data_in <= 24'b000011100001010100101001;
#10000;
	data_in <= 24'b000011000001001100100111;
#10000;
	data_in <= 24'b000100000001010100101010;
#10000;
	data_in <= 24'b000011000001000100100110;
#10000;
	data_in <= 24'b000001110000111100100110;
#10000;
	data_in <= 24'b000100110001101100110010;
#10000;
	data_in <= 24'b000011100001010100101001;
#10000;
	data_in <= 24'b000010000000111100100011;
#10000;
	data_in <= 24'b000011110001011000101001;
#10000;
	data_in <= 24'b000010010001000000100011;
#10000;
	data_in <= 24'b000000110000101000011101;
#10000;
	data_in <= 24'b000011110001011000101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001100000001100010011;
#10000;
	data_in <= 24'b000001000000001100010011;
#10000;
	data_in <= 24'b000001000000010000010110;
#10000;
	data_in <= 24'b000001000000010100011001;
#10000;
	data_in <= 24'b000001010000011000011011;
#10000;
	data_in <= 24'b000001110000011100011111;
#10000;
	data_in <= 24'b000010100000101100100000;
#10000;
	data_in <= 24'b000010110000110100100101;
#10000;
	data_in <= 24'b000001110000011000010110;
#10000;
	data_in <= 24'b000001110000011000010110;
#10000;
	data_in <= 24'b000001100000010100011001;
#10000;
	data_in <= 24'b000001110000011000011010;
#10000;
	data_in <= 24'b000001000000010000011100;
#10000;
	data_in <= 24'b000001000000010000011100;
#10000;
	data_in <= 24'b000000110000010100011101;
#10000;
	data_in <= 24'b000001010000011100011111;
#10000;
	data_in <= 24'b000001100000010100010101;
#10000;
	data_in <= 24'b000001010000010000010100;
#10000;
	data_in <= 24'b000001010000010000011000;
#10000;
	data_in <= 24'b000001110000011000011010;
#10000;
	data_in <= 24'b000001010000010100011101;
#10000;
	data_in <= 24'b000001000000010000011100;
#10000;
	data_in <= 24'b000000110000010000011110;
#10000;
	data_in <= 24'b000001000000010100011111;
#10000;
	data_in <= 24'b000001000000001100010011;
#10000;
	data_in <= 24'b000001000000001000010101;
#10000;
	data_in <= 24'b000001000000001100010111;
#10000;
	data_in <= 24'b000001100000010000011010;
#10000;
	data_in <= 24'b000001100000011000011110;
#10000;
	data_in <= 24'b000001100000010100011111;
#10000;
	data_in <= 24'b000001010000011000100000;
#10000;
	data_in <= 24'b000001110000100000100010;
#10000;
	data_in <= 24'b000001110000011100011001;
#10000;
	data_in <= 24'b000001100000011000011000;
#10000;
	data_in <= 24'b000001010000010000011000;
#10000;
	data_in <= 24'b000001100000010000011010;
#10000;
	data_in <= 24'b000001010000010000011110;
#10000;
	data_in <= 24'b000001100000010000100001;
#10000;
	data_in <= 24'b000001010000011000100010;
#10000;
	data_in <= 24'b000001010000100000100100;
#10000;
	data_in <= 24'b000010000000100000011010;
#10000;
	data_in <= 24'b000001100000010100011001;
#10000;
	data_in <= 24'b000001010000001100011001;
#10000;
	data_in <= 24'b000001000000010000011100;
#10000;
	data_in <= 24'b000001100000010000100001;
#10000;
	data_in <= 24'b000001010000010100100011;
#10000;
	data_in <= 24'b000001000000011000100100;
#10000;
	data_in <= 24'b000001100000100000100110;
#10000;
	data_in <= 24'b000001100000010100011001;
#10000;
	data_in <= 24'b000001000000001100010111;
#10000;
	data_in <= 24'b000000100000001100011000;
#10000;
	data_in <= 24'b000001000000010000011100;
#10000;
	data_in <= 24'b000001100000010000100001;
#10000;
	data_in <= 24'b000001100000011000100100;
#10000;
	data_in <= 24'b000001010000011100100110;
#10000;
	data_in <= 24'b000001100000100000100111;
#10000;
	data_in <= 24'b000001010000010000011000;
#10000;
	data_in <= 24'b000001000000001000011000;
#10000;
	data_in <= 24'b000000100000001000011010;
#10000;
	data_in <= 24'b000001010000010000011110;
#10000;
	data_in <= 24'b000001000000010000100010;
#10000;
	data_in <= 24'b000001010000010000100100;
#10000;
	data_in <= 24'b000000110000010000100110;
#10000;
	data_in <= 24'b000000110000001100100111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001110000101100100100;
#10000;
	data_in <= 24'b000001110000110000100101;
#10000;
	data_in <= 24'b000001110000101100100100;
#10000;
	data_in <= 24'b000001000000011100100011;
#10000;
	data_in <= 24'b000001100000011100100011;
#10000;
	data_in <= 24'b000001100000011000100100;
#10000;
	data_in <= 24'b000010100000110000101011;
#10000;
	data_in <= 24'b000100110001011000110101;
#10000;
	data_in <= 24'b000001100000101000100010;
#10000;
	data_in <= 24'b000010000000110000100100;
#10000;
	data_in <= 24'b000001110000101100100100;
#10000;
	data_in <= 24'b000010000000101100100111;
#10000;
	data_in <= 24'b000010010000101100101001;
#10000;
	data_in <= 24'b000010000000101000101001;
#10000;
	data_in <= 24'b000010010000101000101100;
#10000;
	data_in <= 24'b000011010000111100110001;
#10000;
	data_in <= 24'b000001100000101000100011;
#10000;
	data_in <= 24'b000001110000101100100100;
#10000;
	data_in <= 24'b000001110000101000100110;
#10000;
	data_in <= 24'b000010010000110000101000;
#10000;
	data_in <= 24'b000011000000111000101100;
#10000;
	data_in <= 24'b000010100000110000101011;
#10000;
	data_in <= 24'b000010000000100100101011;
#10000;
	data_in <= 24'b000010000000101000101101;
#10000;
	data_in <= 24'b000001100000100100100101;
#10000;
	data_in <= 24'b000001110000101000100110;
#10000;
	data_in <= 24'b000001100000100100100101;
#10000;
	data_in <= 24'b000001100000100000100110;
#10000;
	data_in <= 24'b000010100000110000101011;
#10000;
	data_in <= 24'b000010100000101100101101;
#10000;
	data_in <= 24'b000010000000100000101100;
#10000;
	data_in <= 24'b000010000000100100101111;
#10000;
	data_in <= 24'b000001010000011100100101;
#10000;
	data_in <= 24'b000001110000100100100111;
#10000;
	data_in <= 24'b000001100000101000100111;
#10000;
	data_in <= 24'b000001100000100100101000;
#10000;
	data_in <= 24'b000010000000101000101100;
#10000;
	data_in <= 24'b000010010000101100101110;
#10000;
	data_in <= 24'b000010010000100100110001;
#10000;
	data_in <= 24'b000010110000101000110100;
#10000;
	data_in <= 24'b000001000000011000100101;
#10000;
	data_in <= 24'b000001110000101000101001;
#10000;
	data_in <= 24'b000010010000110000101011;
#10000;
	data_in <= 24'b000010010000101100101101;
#10000;
	data_in <= 24'b000010110000110100110000;
#10000;
	data_in <= 24'b000010110000110000110010;
#10000;
	data_in <= 24'b000010100000100100110011;
#10000;
	data_in <= 24'b000010100000101100110111;
#10000;
	data_in <= 24'b000001000000011000101000;
#10000;
	data_in <= 24'b000010000000101000101100;
#10000;
	data_in <= 24'b000010010000101100101110;
#10000;
	data_in <= 24'b000001110000101000110000;
#10000;
	data_in <= 24'b000010100000110000110100;
#10000;
	data_in <= 24'b000010100000110000110101;
#10000;
	data_in <= 24'b000010010000100100110111;
#10000;
	data_in <= 24'b000010000000101000111010;
#10000;
	data_in <= 24'b000001100000100000101011;
#10000;
	data_in <= 24'b000010010000101100101110;
#10000;
	data_in <= 24'b000001100000100100101111;
#10000;
	data_in <= 24'b000001010000011100101111;
#10000;
	data_in <= 24'b000010000000101000110011;
#10000;
	data_in <= 24'b000010000000101100111000;
#10000;
	data_in <= 24'b000010000000101000111010;
#10000;
	data_in <= 24'b000001100000101000111011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001110000110000101101;
#10000;
	data_in <= 24'b000001000000100100101010;
#10000;
	data_in <= 24'b000010010001000100101111;
#10000;
	data_in <= 24'b000011010001010100110011;
#10000;
	data_in <= 24'b000010010001000000110001;
#10000;
	data_in <= 24'b000011000001001000110101;
#10000;
	data_in <= 24'b000011100001010000110111;
#10000;
	data_in <= 24'b000010000000111000110001;
#10000;
	data_in <= 24'b000011100001000000110010;
#10000;
	data_in <= 24'b000001010000101000101011;
#10000;
	data_in <= 24'b000000110000100100101100;
#10000;
	data_in <= 24'b000001000000101000101101;
#10000;
	data_in <= 24'b000001110000110100110000;
#10000;
	data_in <= 24'b000100100001101100111101;
#10000;
	data_in <= 24'b000101110001111101000100;
#10000;
	data_in <= 24'b000011000001010100111010;
#10000;
	data_in <= 24'b000101100001100000111011;
#10000;
	data_in <= 24'b000011110001001100110110;
#10000;
	data_in <= 24'b000011010001001100111000;
#10000;
	data_in <= 24'b000010110001000100110110;
#10000;
	data_in <= 24'b000001000000110000110001;
#10000;
	data_in <= 24'b000001110000111100110100;
#10000;
	data_in <= 24'b000011110001011000111101;
#10000;
	data_in <= 24'b000011100001011100111101;
#10000;
	data_in <= 24'b000011100001000000111000;
#10000;
	data_in <= 24'b000010110000110100110101;
#10000;
	data_in <= 24'b000100000001010100111100;
#10000;
	data_in <= 24'b000101110001110001000011;
#10000;
	data_in <= 24'b000010110001000100111010;
#10000;
	data_in <= 24'b000000100000100000110001;
#10000;
	data_in <= 24'b000001110000111000111001;
#10000;
	data_in <= 24'b000100010001101001000101;
#10000;
	data_in <= 24'b000010110000110000111000;
#10000;
	data_in <= 24'b000001000000011100110011;
#10000;
	data_in <= 24'b000010100000110100111001;
#10000;
	data_in <= 24'b000101010001100001000100;
#10000;
	data_in <= 24'b000100100001011101000100;
#10000;
	data_in <= 24'b000010100000111100111100;
#10000;
	data_in <= 24'b000010100001000000111111;
#10000;
	data_in <= 24'b000011110001011101000110;
#10000;
	data_in <= 24'b000011000000111100111100;
#10000;
	data_in <= 24'b000010110000110100111101;
#10000;
	data_in <= 24'b000010110000110100111101;
#10000;
	data_in <= 24'b000010100000111000111110;
#10000;
	data_in <= 24'b000011100001001001000011;
#10000;
	data_in <= 24'b000011110001010001000101;
#10000;
	data_in <= 24'b000011010001010001000110;
#10000;
	data_in <= 24'b000010100001001001000111;
#10000;
	data_in <= 24'b000001110000100000111010;
#10000;
	data_in <= 24'b000010110000111101000000;
#10000;
	data_in <= 24'b000011000001000001000001;
#10000;
	data_in <= 24'b000010010000110000111111;
#10000;
	data_in <= 24'b000010110000111101000100;
#10000;
	data_in <= 24'b000011110001010101001010;
#10000;
	data_in <= 24'b000100010001011001001101;
#10000;
	data_in <= 24'b000100000001011101010000;
#10000;
	data_in <= 24'b000010010000110000111111;
#10000;
	data_in <= 24'b000011010000111101000101;
#10000;
	data_in <= 24'b000011100001000001000110;
#10000;
	data_in <= 24'b000011100001001001000111;
#10000;
	data_in <= 24'b000011100001001101001010;
#10000;
	data_in <= 24'b000011000001001101001100;
#10000;
	data_in <= 24'b000011000001001001001101;
#10000;
	data_in <= 24'b000011000001010001010000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001100000111100110001;
#10000;
	data_in <= 24'b000010100001001000110111;
#10000;
	data_in <= 24'b000100000001100000111101;
#10000;
	data_in <= 24'b000101000001110101000011;
#10000;
	data_in <= 24'b000100110001110101000101;
#10000;
	data_in <= 24'b000101000001110101001000;
#10000;
	data_in <= 24'b000101000001111001001101;
#10000;
	data_in <= 24'b000101110010000101010001;
#10000;
	data_in <= 24'b000010110001010000111010;
#10000;
	data_in <= 24'b000011000001010100111011;
#10000;
	data_in <= 24'b000011100001011000111110;
#10000;
	data_in <= 24'b000011100001011101000010;
#10000;
	data_in <= 24'b000011100001011101000011;
#10000;
	data_in <= 24'b000011010001010101000100;
#10000;
	data_in <= 24'b000011110001011001000111;
#10000;
	data_in <= 24'b000011110001100101001001;
#10000;
	data_in <= 24'b000010010001000100111001;
#10000;
	data_in <= 24'b000001010000111000111001;
#10000;
	data_in <= 24'b000001010000111000111010;
#10000;
	data_in <= 24'b000001010000111100111110;
#10000;
	data_in <= 24'b000001110001000101000001;
#10000;
	data_in <= 24'b000010010001001101000011;
#10000;
	data_in <= 24'b000010110001010001000110;
#10000;
	data_in <= 24'b000011000001011101001001;
#10000;
	data_in <= 24'b000100010001101001000110;
#10000;
	data_in <= 24'b000011000001011001000101;
#10000;
	data_in <= 24'b000010100001010001000100;
#10000;
	data_in <= 24'b000010100001001101000101;
#10000;
	data_in <= 24'b000011000001010001001001;
#10000;
	data_in <= 24'b000010110001011001001010;
#10000;
	data_in <= 24'b000011000001011001001100;
#10000;
	data_in <= 24'b000011000001100001001110;
#10000;
	data_in <= 24'b000100100001100101001010;
#10000;
	data_in <= 24'b000011100001011101001001;
#10000;
	data_in <= 24'b000011010001010101001010;
#10000;
	data_in <= 24'b000011000001011001001100;
#10000;
	data_in <= 24'b000011110001100001010001;
#10000;
	data_in <= 24'b000011100001100101010011;
#10000;
	data_in <= 24'b000100000001101001010110;
#10000;
	data_in <= 24'b000100000001101101010111;
#10000;
	data_in <= 24'b000011010001010001001011;
#10000;
	data_in <= 24'b000010100001001101001100;
#10000;
	data_in <= 24'b000010110001001101001110;
#10000;
	data_in <= 24'b000011000001011001010010;
#10000;
	data_in <= 24'b000100000001100101011000;
#10000;
	data_in <= 24'b000100100001110101011011;
#10000;
	data_in <= 24'b000101000001111001011110;
#10000;
	data_in <= 24'b000100110001111101011111;
#10000;
	data_in <= 24'b000101000001110001010111;
#10000;
	data_in <= 24'b000100010001101101010111;
#10000;
	data_in <= 24'b000011110001101001011000;
#10000;
	data_in <= 24'b000011110001101101011011;
#10000;
	data_in <= 24'b000011110001101101011101;
#10000;
	data_in <= 24'b000011110001101101011101;
#10000;
	data_in <= 24'b000100000001101101011111;
#10000;
	data_in <= 24'b000100000001110001100010;
#10000;
	data_in <= 24'b000011010001011001010110;
#10000;
	data_in <= 24'b000010110001010101010101;
#10000;
	data_in <= 24'b000010010001010001011000;
#10000;
	data_in <= 24'b000010010001011001011010;
#10000;
	data_in <= 24'b000010010001010101011011;
#10000;
	data_in <= 24'b000010000001011101011100;
#10000;
	data_in <= 24'b000010100001100001100000;
#10000;
	data_in <= 24'b000011000001100101100011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000100010001111101001111;
#10000;
	data_in <= 24'b000100000001111101010000;
#10000;
	data_in <= 24'b000100010010000001010001;
#10000;
	data_in <= 24'b000100110010010001010111;
#10000;
	data_in <= 24'b000101010010010101011010;
#10000;
	data_in <= 24'b000101010010011001011110;
#10000;
	data_in <= 24'b000101110010100101100100;
#10000;
	data_in <= 24'b000110000010111001101000;
#10000;
	data_in <= 24'b000101000001111101010001;
#10000;
	data_in <= 24'b000100000001111001001111;
#10000;
	data_in <= 24'b000011100001110001010000;
#10000;
	data_in <= 24'b000011010001110101010010;
#10000;
	data_in <= 24'b000011110010000001011000;
#10000;
	data_in <= 24'b000100010010010001011101;
#10000;
	data_in <= 24'b000110000010101101101000;
#10000;
	data_in <= 24'b000110100011000101101111;
#10000;
	data_in <= 24'b000011000001011101001011;
#10000;
	data_in <= 24'b000010110001011101001101;
#10000;
	data_in <= 24'b000010110001100101001110;
#10000;
	data_in <= 24'b000011000001101101010011;
#10000;
	data_in <= 24'b000011000001110101010110;
#10000;
	data_in <= 24'b000010110001110101011000;
#10000;
	data_in <= 24'b000011010010000001011101;
#10000;
	data_in <= 24'b000011000010001101100001;
#10000;
	data_in <= 24'b000011000001011101010000;
#10000;
	data_in <= 24'b000011100001101101010011;
#10000;
	data_in <= 24'b000100000001111001011000;
#10000;
	data_in <= 24'b000100010010000101011100;
#10000;
	data_in <= 24'b000100000010001001011111;
#10000;
	data_in <= 24'b000011100010000101011110;
#10000;
	data_in <= 24'b000011000010000001100001;
#10000;
	data_in <= 24'b000010010001111101100000;
#10000;
	data_in <= 24'b000100010001111001011100;
#10000;
	data_in <= 24'b000100000001111101011101;
#10000;
	data_in <= 24'b000100010010000001011111;
#10000;
	data_in <= 24'b000100000010000101100000;
#10000;
	data_in <= 24'b000100010010001101100100;
#10000;
	data_in <= 24'b000100100010011001100111;
#10000;
	data_in <= 24'b000101010010100001101100;
#10000;
	data_in <= 24'b000101000010100101101101;
#10000;
	data_in <= 24'b000100010001111101100001;
#10000;
	data_in <= 24'b000100000010000001100011;
#10000;
	data_in <= 24'b000100000010000001100011;
#10000;
	data_in <= 24'b000011110001111101100100;
#10000;
	data_in <= 24'b000011100010000101100101;
#10000;
	data_in <= 24'b000100000010010001101011;
#10000;
	data_in <= 24'b000100110010011001101111;
#10000;
	data_in <= 24'b000100100010100001110000;
#10000;
	data_in <= 24'b000011110001111001100110;
#10000;
	data_in <= 24'b000100010010000001101001;
#10000;
	data_in <= 24'b000101000010001101101100;
#10000;
	data_in <= 24'b000100100010001001101110;
#10000;
	data_in <= 24'b000100110010001101101111;
#10000;
	data_in <= 24'b000100100010010001110001;
#10000;
	data_in <= 24'b000100110010010101110010;
#10000;
	data_in <= 24'b000100000010010001110001;
#10000;
	data_in <= 24'b000010010001100101100110;
#10000;
	data_in <= 24'b000010100001101101101010;
#10000;
	data_in <= 24'b000011110001111001101101;
#10000;
	data_in <= 24'b000011100001111101110000;
#10000;
	data_in <= 24'b000011110010000001110001;
#10000;
	data_in <= 24'b000100000010001101110100;
#10000;
	data_in <= 24'b000100100010010101110110;
#10000;
	data_in <= 24'b000100010010001101110110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000101110011000101101101;
#10000;
	data_in <= 24'b000110100011011001110010;
#10000;
	data_in <= 24'b000101010011000101101110;
#10000;
	data_in <= 24'b000110100011010101110101;
#10000;
	data_in <= 24'b001001100100000110000001;
#10000;
	data_in <= 24'b000111100011100001111010;
#10000;
	data_in <= 24'b000100100010111001101110;
#10000;
	data_in <= 24'b000110010011011001110011;
#10000;
	data_in <= 24'b000110000010111101101101;
#10000;
	data_in <= 24'b000110110011010001110100;
#10000;
	data_in <= 24'b000110100011001101110011;
#10000;
	data_in <= 24'b000111100011011101110111;
#10000;
	data_in <= 24'b001000110011110001111100;
#10000;
	data_in <= 24'b000110000011000101110001;
#10000;
	data_in <= 24'b000011010010011001100110;
#10000;
	data_in <= 24'b000101000010101101101001;
#10000;
	data_in <= 24'b000011110010010101100110;
#10000;
	data_in <= 24'b000011010010010101100111;
#10000;
	data_in <= 24'b000011000010010001100110;
#10000;
	data_in <= 24'b000100000010100001101010;
#10000;
	data_in <= 24'b000100110010101101101101;
#10000;
	data_in <= 24'b000011110010100001101000;
#10000;
	data_in <= 24'b000010110010010001100100;
#10000;
	data_in <= 24'b000011110010011001100100;
#10000;
	data_in <= 24'b000100010010100101101011;
#10000;
	data_in <= 24'b000010110010001001100110;
#10000;
	data_in <= 24'b000010000001111101100011;
#10000;
	data_in <= 24'b000010100010000101100101;
#10000;
	data_in <= 24'b000011010010010001101000;
#10000;
	data_in <= 24'b000011100010011001101000;
#10000;
	data_in <= 24'b000011000010010001100110;
#10000;
	data_in <= 24'b000011000010001001100100;
#10000;
	data_in <= 24'b000100110010100101110000;
#10000;
	data_in <= 24'b000100000010011001101101;
#10000;
	data_in <= 24'b000100100010100001101111;
#10000;
	data_in <= 24'b000101010010101101110010;
#10000;
	data_in <= 24'b000101010010101101110010;
#10000;
	data_in <= 24'b000101100010110101110001;
#10000;
	data_in <= 24'b000101010010110001110000;
#10000;
	data_in <= 24'b000100110010100001101100;
#10000;
	data_in <= 24'b000011100010001101101110;
#10000;
	data_in <= 24'b000100000010010101110000;
#10000;
	data_in <= 24'b000101000010100101110100;
#10000;
	data_in <= 24'b000101000010100101110100;
#10000;
	data_in <= 24'b000100010010011101101111;
#10000;
	data_in <= 24'b000100100010100001110000;
#10000;
	data_in <= 24'b000101100010110001110100;
#10000;
	data_in <= 24'b000101100010110001110100;
#10000;
	data_in <= 24'b000100100010011001110100;
#10000;
	data_in <= 24'b000100100010100001110110;
#10000;
	data_in <= 24'b000100000010011001110100;
#10000;
	data_in <= 24'b000011000010001001110000;
#10000;
	data_in <= 24'b000010110001111101101100;
#10000;
	data_in <= 24'b000011000010000001101101;
#10000;
	data_in <= 24'b000011010010000101101110;
#10000;
	data_in <= 24'b000011100010001001101111;
#10000;
	data_in <= 24'b000100010010011001111000;
#10000;
	data_in <= 24'b000100100010011101111001;
#10000;
	data_in <= 24'b000100000010010101110111;
#10000;
	data_in <= 24'b000100000010010101110111;
#10000;
	data_in <= 24'b000101100010100001111011;
#10000;
	data_in <= 24'b000101110010101001111011;
#10000;
	data_in <= 24'b000100100010010101110110;
#10000;
	data_in <= 24'b000011010010000001110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000101100011000001101100;
#10000;
	data_in <= 24'b000101100010110001100110;
#10000;
	data_in <= 24'b000100110010011001011111;
#10000;
	data_in <= 24'b000101000010001101011011;
#10000;
	data_in <= 24'b000101000010010001011001;
#10000;
	data_in <= 24'b000100110010010001010111;
#10000;
	data_in <= 24'b000100110010001001010011;
#10000;
	data_in <= 24'b000100010010000101010000;
#10000;
	data_in <= 24'b000110010010110101100111;
#10000;
	data_in <= 24'b000110010010110001100101;
#10000;
	data_in <= 24'b000101110010100001100001;
#10000;
	data_in <= 24'b000100100010001101011011;
#10000;
	data_in <= 24'b000100110010001101011000;
#10000;
	data_in <= 24'b000101000010010101011000;
#10000;
	data_in <= 24'b000101010010001101010111;
#10000;
	data_in <= 24'b000100110010001001010011;
#10000;
	data_in <= 24'b000011100010001101100001;
#10000;
	data_in <= 24'b000100010010010001100001;
#10000;
	data_in <= 24'b000100000010001001011111;
#10000;
	data_in <= 24'b000011000001111001011001;
#10000;
	data_in <= 24'b000011000001110101010110;
#10000;
	data_in <= 24'b000100000001111101010111;
#10000;
	data_in <= 24'b000100100010000001010101;
#10000;
	data_in <= 24'b000100010001111101010011;
#10000;
	data_in <= 24'b000011000010000001100001;
#10000;
	data_in <= 24'b000011010001111101100000;
#10000;
	data_in <= 24'b000011010001111001011101;
#10000;
	data_in <= 24'b000011010001111001011101;
#10000;
	data_in <= 24'b000011110001111001011100;
#10000;
	data_in <= 24'b000011010001110101011000;
#10000;
	data_in <= 24'b000011100001110001010110;
#10000;
	data_in <= 24'b000100000001110101010101;
#10000;
	data_in <= 24'b000101100010100101101101;
#10000;
	data_in <= 24'b000100000010001101100111;
#10000;
	data_in <= 24'b000100010010001001100101;
#10000;
	data_in <= 24'b000101100010011101101010;
#10000;
	data_in <= 24'b000101110010011101101001;
#10000;
	data_in <= 24'b000100100010000101100000;
#10000;
	data_in <= 24'b000011110001110001011010;
#10000;
	data_in <= 24'b000100100001110101011001;
#10000;
	data_in <= 24'b000101110010101001110011;
#10000;
	data_in <= 24'b000100100010001101101100;
#10000;
	data_in <= 24'b000100110010001001101010;
#10000;
	data_in <= 24'b000110000010011101101111;
#10000;
	data_in <= 24'b000110000010011101101100;
#10000;
	data_in <= 24'b000011110001111101100010;
#10000;
	data_in <= 24'b000010100001011101011011;
#10000;
	data_in <= 24'b000011000001100001011000;
#10000;
	data_in <= 24'b000100010010001101110000;
#10000;
	data_in <= 24'b000011100010000001101101;
#10000;
	data_in <= 24'b000011110001111101101011;
#10000;
	data_in <= 24'b000100010010000101101101;
#10000;
	data_in <= 24'b000100010010000001101001;
#10000;
	data_in <= 24'b000011000001101001100010;
#10000;
	data_in <= 24'b000010010001010101011101;
#10000;
	data_in <= 24'b000010010001010001011000;
#10000;
	data_in <= 24'b000011100001111101110000;
#10000;
	data_in <= 24'b000100000010000101110010;
#10000;
	data_in <= 24'b000100000010000101110010;
#10000;
	data_in <= 24'b000100000001111101101110;
#10000;
	data_in <= 24'b000011100001111001101011;
#10000;
	data_in <= 24'b000011110001110101101001;
#10000;
	data_in <= 24'b000011010001101001100110;
#10000;
	data_in <= 24'b000010110001011101011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000011110001111001001100;
#10000;
	data_in <= 24'b000101000010000101001101;
#10000;
	data_in <= 24'b000101110010001101001101;
#10000;
	data_in <= 24'b000101000001111001000110;
#10000;
	data_in <= 24'b000010110001011000111100;
#10000;
	data_in <= 24'b000001110001001000111000;
#10000;
	data_in <= 24'b000010000001010000111000;
#10000;
	data_in <= 24'b000011100001011100111100;
#10000;
	data_in <= 24'b000110010010010101010101;
#10000;
	data_in <= 24'b000100100001111101001101;
#10000;
	data_in <= 24'b000011010001100001000100;
#10000;
	data_in <= 24'b000011000001010101000000;
#10000;
	data_in <= 24'b000011100001011000111110;
#10000;
	data_in <= 24'b000011100001011000111110;
#10000;
	data_in <= 24'b000011000001010000111100;
#10000;
	data_in <= 24'b000010100001001100111001;
#10000;
	data_in <= 24'b000011110001101001001100;
#10000;
	data_in <= 24'b000011010001100101001001;
#10000;
	data_in <= 24'b000011010001011101000111;
#10000;
	data_in <= 24'b000011100001011001000101;
#10000;
	data_in <= 24'b000100000001011001000011;
#10000;
	data_in <= 24'b000011110001011001000001;
#10000;
	data_in <= 24'b000011100001010101000000;
#10000;
	data_in <= 24'b000011000001010000111100;
#10000;
	data_in <= 24'b000010000001010001001010;
#10000;
	data_in <= 24'b000011100001100101001101;
#10000;
	data_in <= 24'b000100110001110001001110;
#10000;
	data_in <= 24'b000100100001110001001100;
#10000;
	data_in <= 24'b000100000001011101001000;
#10000;
	data_in <= 24'b000011110001010101000100;
#10000;
	data_in <= 24'b000100000001011001000011;
#10000;
	data_in <= 24'b000100100001100001000101;
#10000;
	data_in <= 24'b000100110001111001011000;
#10000;
	data_in <= 24'b000100100001101101010100;
#10000;
	data_in <= 24'b000100000001011101001110;
#10000;
	data_in <= 24'b000011010001010101001010;
#10000;
	data_in <= 24'b000011110001010101001010;
#10000;
	data_in <= 24'b000100000001011101001001;
#10000;
	data_in <= 24'b000100010001011001000111;
#10000;
	data_in <= 24'b000100000001010101000110;
#10000;
	data_in <= 24'b000011110001101001011000;
#10000;
	data_in <= 24'b000011000001011001010010;
#10000;
	data_in <= 24'b000010010001000101001100;
#10000;
	data_in <= 24'b000010110001001001001011;
#10000;
	data_in <= 24'b000011100001001101001010;
#10000;
	data_in <= 24'b000011110001010001001011;
#10000;
	data_in <= 24'b000011110001001101001000;
#10000;
	data_in <= 24'b000011000001000001000011;
#10000;
	data_in <= 24'b000001100000111101010010;
#10000;
	data_in <= 24'b000010000001000101010001;
#10000;
	data_in <= 24'b000010110001001001010001;
#10000;
	data_in <= 24'b000010110001001101001111;
#10000;
	data_in <= 24'b000011000001001001001101;
#10000;
	data_in <= 24'b000010110001000101001100;
#10000;
	data_in <= 24'b000011010001000101001011;
#10000;
	data_in <= 24'b000011010001001001001001;
#10000;
	data_in <= 24'b000011000001011001011100;
#10000;
	data_in <= 24'b000011000001010101011001;
#10000;
	data_in <= 24'b000010110001001101010110;
#10000;
	data_in <= 24'b000010100001000001010001;
#10000;
	data_in <= 24'b000010010001000001001111;
#10000;
	data_in <= 24'b000011000001000101010000;
#10000;
	data_in <= 24'b000011110001010001010001;
#10000;
	data_in <= 24'b000100000001011001010001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000100010001011100111010;
#10000;
	data_in <= 24'b000011010001001100110110;
#10000;
	data_in <= 24'b000010110001001000110011;
#10000;
	data_in <= 24'b000011010001010000110101;
#10000;
	data_in <= 24'b000011100001010100110110;
#10000;
	data_in <= 24'b000011010001010100110011;
#10000;
	data_in <= 24'b000011000001010000110010;
#10000;
	data_in <= 24'b000011010001010100110010;
#10000;
	data_in <= 24'b000010010001000100110110;
#10000;
	data_in <= 24'b000010000001000100110011;
#10000;
	data_in <= 24'b000010100001001100110101;
#10000;
	data_in <= 24'b000011100001011100111000;
#10000;
	data_in <= 24'b000100010001100000111001;
#10000;
	data_in <= 24'b000011010001010100110011;
#10000;
	data_in <= 24'b000010010001000100101111;
#10000;
	data_in <= 24'b000010000001000000101101;
#10000;
	data_in <= 24'b000011100001010000111101;
#10000;
	data_in <= 24'b000011000001001100111010;
#10000;
	data_in <= 24'b000011000001001100111010;
#10000;
	data_in <= 24'b000011100001011000111011;
#10000;
	data_in <= 24'b000011100001011100111001;
#10000;
	data_in <= 24'b000010110001010000110101;
#10000;
	data_in <= 24'b000010100001000100110010;
#10000;
	data_in <= 24'b000010010001000100101111;
#10000;
	data_in <= 24'b000100010001011101000010;
#10000;
	data_in <= 24'b000011100001010000111101;
#10000;
	data_in <= 24'b000011010001001100111100;
#10000;
	data_in <= 24'b000011000001001100111010;
#10000;
	data_in <= 24'b000010110001001100111000;
#10000;
	data_in <= 24'b000010010001000100110110;
#10000;
	data_in <= 24'b000010010000111100110010;
#10000;
	data_in <= 24'b000010000000111100110000;
#10000;
	data_in <= 24'b000010110001000101000000;
#10000;
	data_in <= 24'b000010100001000000111101;
#10000;
	data_in <= 24'b000010100001000000111101;
#10000;
	data_in <= 24'b000010110001001000111101;
#10000;
	data_in <= 24'b000010110001000100111010;
#10000;
	data_in <= 24'b000001110000110100110110;
#10000;
	data_in <= 24'b000001100000101100110010;
#10000;
	data_in <= 24'b000001010000101100110000;
#10000;
	data_in <= 24'b000011100001001001000101;
#10000;
	data_in <= 24'b000011010001001001000011;
#10000;
	data_in <= 24'b000011000001001001000001;
#10000;
	data_in <= 24'b000010110001000101000000;
#10000;
	data_in <= 24'b000010110001000000111101;
#10000;
	data_in <= 24'b000010110001000100111100;
#10000;
	data_in <= 24'b000011010001000100111010;
#10000;
	data_in <= 24'b000011010001001000111001;
#10000;
	data_in <= 24'b000100100001011101001110;
#10000;
	data_in <= 24'b000100000001011001001011;
#10000;
	data_in <= 24'b000011010001010001000110;
#10000;
	data_in <= 24'b000010100001000101000011;
#10000;
	data_in <= 24'b000011000001000101000010;
#10000;
	data_in <= 24'b000011010001001101000010;
#10000;
	data_in <= 24'b000100010001011101000010;
#10000;
	data_in <= 24'b000100100001100001000001;
#10000;
	data_in <= 24'b000011010001010001001101;
#10000;
	data_in <= 24'b000011010001010001001011;
#10000;
	data_in <= 24'b000011010001010001001011;
#10000;
	data_in <= 24'b000011010001001101001000;
#10000;
	data_in <= 24'b000011000001001101000101;
#10000;
	data_in <= 24'b000011010001001001000011;
#10000;
	data_in <= 24'b000011010001000101000001;
#10000;
	data_in <= 24'b000011010001001100111110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000100000001100100110100;
#10000;
	data_in <= 24'b000100000001100100110100;
#10000;
	data_in <= 24'b000100000001011100110010;
#10000;
	data_in <= 24'b000011110001011000110001;
#10000;
	data_in <= 24'b000011000001001100101110;
#10000;
	data_in <= 24'b000010110001000000101001;
#10000;
	data_in <= 24'b000010010000111000100111;
#10000;
	data_in <= 24'b000010010000110100100101;
#10000;
	data_in <= 24'b000011010001010000101111;
#10000;
	data_in <= 24'b000010110001001000101101;
#10000;
	data_in <= 24'b000010110001001000101101;
#10000;
	data_in <= 24'b000010110001001000101011;
#10000;
	data_in <= 24'b000011000001000100101010;
#10000;
	data_in <= 24'b000010100000111100101000;
#10000;
	data_in <= 24'b000010100000111000100111;
#10000;
	data_in <= 24'b000010110000111100100111;
#10000;
	data_in <= 24'b000010110001000000101111;
#10000;
	data_in <= 24'b000010000000111000101011;
#10000;
	data_in <= 24'b000010010000110100101010;
#10000;
	data_in <= 24'b000011000001000000101100;
#10000;
	data_in <= 24'b000011000001000000101100;
#10000;
	data_in <= 24'b000010010000110100101001;
#10000;
	data_in <= 24'b000010100000110100101001;
#10000;
	data_in <= 24'b000011000001000000101001;
#10000;
	data_in <= 24'b000011100001001100110100;
#10000;
	data_in <= 24'b000010010000111000101101;
#10000;
	data_in <= 24'b000010100000110100101100;
#10000;
	data_in <= 24'b000011000001000000101101;
#10000;
	data_in <= 24'b000010110000111100101100;
#10000;
	data_in <= 24'b000001110000101100100111;
#10000;
	data_in <= 24'b000010000000101000101000;
#10000;
	data_in <= 24'b000010110000111000101010;
#10000;
	data_in <= 24'b000100010001010100111000;
#10000;
	data_in <= 24'b000011010001001000110011;
#10000;
	data_in <= 24'b000011000000111000110000;
#10000;
	data_in <= 24'b000011010001000000101111;
#10000;
	data_in <= 24'b000010110000111000101101;
#10000;
	data_in <= 24'b000001110000101100101000;
#10000;
	data_in <= 24'b000001100000100100101000;
#10000;
	data_in <= 24'b000001110000101100101000;
#10000;
	data_in <= 24'b000100110001011000111100;
#10000;
	data_in <= 24'b000100000001010000110111;
#10000;
	data_in <= 24'b000011110001000100110100;
#10000;
	data_in <= 24'b000011100001000000110010;
#10000;
	data_in <= 24'b000011010000111100110001;
#10000;
	data_in <= 24'b000010110000111000101101;
#10000;
	data_in <= 24'b000010010000110000101011;
#10000;
	data_in <= 24'b000010000000101100101010;
#10000;
	data_in <= 24'b000011100001001100111010;
#10000;
	data_in <= 24'b000011100001010000111001;
#10000;
	data_in <= 24'b000011100001000100110111;
#10000;
	data_in <= 24'b000011000001000000110011;
#10000;
	data_in <= 24'b000011010000111100110010;
#10000;
	data_in <= 24'b000011010000111100110001;
#10000;
	data_in <= 24'b000010110000110100101111;
#10000;
	data_in <= 24'b000010000000101100101010;
#10000;
	data_in <= 24'b000010100000111000110111;
#10000;
	data_in <= 24'b000010110001000000110111;
#10000;
	data_in <= 24'b000010110000110100110101;
#10000;
	data_in <= 24'b000010000000101100110001;
#10000;
	data_in <= 24'b000010100000101100110001;
#10000;
	data_in <= 24'b000011000000111000110001;
#10000;
	data_in <= 24'b000010010000101100101110;
#10000;
	data_in <= 24'b000001000000011000101000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000100000001010100101010;
#10000;
	data_in <= 24'b000011110001001000100111;
#10000;
	data_in <= 24'b000010100000110100100010;
#10000;
	data_in <= 24'b000001010000101000011111;
#10000;
	data_in <= 24'b000000110000100000011101;
#10000;
	data_in <= 24'b000001000000100100011110;
#10000;
	data_in <= 24'b000001110000110000100001;
#10000;
	data_in <= 24'b000010010000111000100011;
#10000;
	data_in <= 24'b000011000000111000100110;
#10000;
	data_in <= 24'b000011000000111100100100;
#10000;
	data_in <= 24'b000010110000111000100011;
#10000;
	data_in <= 24'b000011000000111100100100;
#10000;
	data_in <= 24'b000011010001000000100101;
#10000;
	data_in <= 24'b000011010001000000100101;
#10000;
	data_in <= 24'b000010110000111000100011;
#10000;
	data_in <= 24'b000010010000110000100001;
#10000;
	data_in <= 24'b000011000000111000100110;
#10000;
	data_in <= 24'b000010010000101100100011;
#10000;
	data_in <= 24'b000010000000101000100010;
#10000;
	data_in <= 24'b000010010000101100100011;
#10000;
	data_in <= 24'b000010110000110100100101;
#10000;
	data_in <= 24'b000011000000111000100110;
#10000;
	data_in <= 24'b000010100000110100100010;
#10000;
	data_in <= 24'b000010000000101100100000;
#10000;
	data_in <= 24'b000010100000101100100101;
#10000;
	data_in <= 24'b000001110000100100100001;
#10000;
	data_in <= 24'b000001010000011100011111;
#10000;
	data_in <= 24'b000001010000011100011111;
#10000;
	data_in <= 24'b000001110000100100100001;
#10000;
	data_in <= 24'b000010010000101100100011;
#10000;
	data_in <= 24'b000010100000110000100100;
#10000;
	data_in <= 24'b000010010000110000100001;
#10000;
	data_in <= 24'b000001100000101000100011;
#10000;
	data_in <= 24'b000001100000101000100011;
#10000;
	data_in <= 24'b000001100000101000100011;
#10000;
	data_in <= 24'b000001110000101100100100;
#10000;
	data_in <= 24'b000010000000110000100101;
#10000;
	data_in <= 24'b000010100000111000100110;
#10000;
	data_in <= 24'b000010100000111000100110;
#10000;
	data_in <= 24'b000010100000111000100110;
#10000;
	data_in <= 24'b000011010001000000101100;
#10000;
	data_in <= 24'b000011000001000000101001;
#10000;
	data_in <= 24'b000010100000110100101001;
#10000;
	data_in <= 24'b000010010000110100100110;
#10000;
	data_in <= 24'b000010000000110000100101;
#10000;
	data_in <= 24'b000010010000110100100110;
#10000;
	data_in <= 24'b000010110000111100101000;
#10000;
	data_in <= 24'b000011000001000000101000;
#10000;
	data_in <= 24'b000011110001001100110000;
#10000;
	data_in <= 24'b000011000001000000101100;
#10000;
	data_in <= 24'b000010010000110100101010;
#10000;
	data_in <= 24'b000001110000101100100111;
#10000;
	data_in <= 24'b000001110000101100100111;
#10000;
	data_in <= 24'b000010010000110100101001;
#10000;
	data_in <= 24'b000010110000111000101010;
#10000;
	data_in <= 24'b000011000001000000101001;
#10000;
	data_in <= 24'b000001100000100100101000;
#10000;
	data_in <= 24'b000001100000100100101000;
#10000;
	data_in <= 24'b000001110000101000101001;
#10000;
	data_in <= 24'b000010100000111000101011;
#10000;
	data_in <= 24'b000011100001001000101111;
#10000;
	data_in <= 24'b000011110001001100110000;
#10000;
	data_in <= 24'b000011010000111100101101;
#10000;
	data_in <= 24'b000010100000110100101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000011000001000100100110;
#10000;
	data_in <= 24'b000010100000111100100100;
#10000;
	data_in <= 24'b000001100000101100100000;
#10000;
	data_in <= 24'b000011100001001100101000;
#10000;
	data_in <= 24'b000011100001001100101000;
#10000;
	data_in <= 24'b000010100000111100100100;
#10000;
	data_in <= 24'b000011100001001100101000;
#10000;
	data_in <= 24'b000010000000110100100010;
#10000;
	data_in <= 24'b000010000000101100100000;
#10000;
	data_in <= 24'b000010010000110000100001;
#10000;
	data_in <= 24'b000010100000110100100010;
#10000;
	data_in <= 24'b000011110001001000100111;
#10000;
	data_in <= 24'b000011010001000000100101;
#10000;
	data_in <= 24'b000010100000110100100010;
#10000;
	data_in <= 24'b000010110000111000100011;
#10000;
	data_in <= 24'b000010010000110000100001;
#10000;
	data_in <= 24'b000010100000110100100010;
#10000;
	data_in <= 24'b000010100000110100100010;
#10000;
	data_in <= 24'b000100000001001100101000;
#10000;
	data_in <= 24'b000011010001000000100101;
#10000;
	data_in <= 24'b000001110000101000011111;
#10000;
	data_in <= 24'b000001110000101000011111;
#10000;
	data_in <= 24'b000001100000100100011110;
#10000;
	data_in <= 24'b000001100000100100011110;
#10000;
	data_in <= 24'b000011100001000100100110;
#10000;
	data_in <= 24'b000010110000111000100011;
#10000;
	data_in <= 24'b000011110001001000100111;
#10000;
	data_in <= 24'b000010000000101100100000;
#10000;
	data_in <= 24'b000000110000011000011011;
#10000;
	data_in <= 24'b000010000000101100100000;
#10000;
	data_in <= 24'b000001010000100000011101;
#10000;
	data_in <= 24'b000001100000100100011110;
#10000;
	data_in <= 24'b000011010000111100100111;
#10000;
	data_in <= 24'b000001100000100000100000;
#10000;
	data_in <= 24'b000010010000101100100011;
#10000;
	data_in <= 24'b000001000000011000011110;
#10000;
	data_in <= 24'b000001000000011100011100;
#10000;
	data_in <= 24'b000010110000111000100011;
#10000;
	data_in <= 24'b000001110000101000011111;
#10000;
	data_in <= 24'b000001010000100000011101;
#10000;
	data_in <= 24'b000011010000111100100111;
#10000;
	data_in <= 24'b000001110000100100100001;
#10000;
	data_in <= 24'b000010000000101000100010;
#10000;
	data_in <= 24'b000001110000100100100001;
#10000;
	data_in <= 24'b000010000000101000100010;
#10000;
	data_in <= 24'b000011000000111100100100;
#10000;
	data_in <= 24'b000001110000101000011111;
#10000;
	data_in <= 24'b000000100000010100011010;
#10000;
	data_in <= 24'b000011010001000100101010;
#10000;
	data_in <= 24'b000010100000111000100111;
#10000;
	data_in <= 24'b000001110000101100100100;
#10000;
	data_in <= 24'b000010010000110100100101;
#10000;
	data_in <= 24'b000010010000101100100011;
#10000;
	data_in <= 24'b000001100000100000100000;
#10000;
	data_in <= 24'b000001100000100000100000;
#10000;
	data_in <= 24'b000000010000001100011011;
#10000;
	data_in <= 24'b000010100000110100101001;
#10000;
	data_in <= 24'b000010100000110100101001;
#10000;
	data_in <= 24'b000001010000100000100100;
#10000;
	data_in <= 24'b000010000000110000100101;
#10000;
	data_in <= 24'b000001100000011100100001;
#10000;
	data_in <= 24'b000000000000001000011010;
#10000;
	data_in <= 24'b000001100000011100100001;
#10000;
	data_in <= 24'b000001000000011000011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001000000001000011000;
#10000;
	data_in <= 24'b000001010000001100011001;
#10000;
	data_in <= 24'b000001000000001100011101;
#10000;
	data_in <= 24'b000001010000001100100000;
#10000;
	data_in <= 24'b000001010000010000100100;
#10000;
	data_in <= 24'b000001100000010100100111;
#10000;
	data_in <= 24'b000001000000010000101000;
#10000;
	data_in <= 24'b000001000000001100101010;
#10000;
	data_in <= 24'b000001100000010000011010;
#10000;
	data_in <= 24'b000001100000001100011100;
#10000;
	data_in <= 24'b000001010000001100100000;
#10000;
	data_in <= 24'b000001100000010000100010;
#10000;
	data_in <= 24'b000001010000010000100110;
#10000;
	data_in <= 24'b000001100000010000101000;
#10000;
	data_in <= 24'b000001010000010000101011;
#10000;
	data_in <= 24'b000001010000010000101100;
#10000;
	data_in <= 24'b000001000000010000011100;
#10000;
	data_in <= 24'b000001000000010000011100;
#10000;
	data_in <= 24'b000001010000001100100000;
#10000;
	data_in <= 24'b000001010000001100100001;
#10000;
	data_in <= 24'b000001000000001100100101;
#10000;
	data_in <= 24'b000001100000010000101000;
#10000;
	data_in <= 24'b000001010000010000101011;
#10000;
	data_in <= 24'b000001100000010100101101;
#10000;
	data_in <= 24'b000000110000001100011011;
#10000;
	data_in <= 24'b000001000000001100011101;
#10000;
	data_in <= 24'b000001000000001000100000;
#10000;
	data_in <= 24'b000001010000001000100010;
#10000;
	data_in <= 24'b000001000000001000100110;
#10000;
	data_in <= 24'b000001010000001000101001;
#10000;
	data_in <= 24'b000001010000010000101100;
#10000;
	data_in <= 24'b000001100000010100101111;
#10000;
	data_in <= 24'b000000110000001000011100;
#10000;
	data_in <= 24'b000001000000001100011101;
#10000;
	data_in <= 24'b000001010000001100100001;
#10000;
	data_in <= 24'b000001010000001000100010;
#10000;
	data_in <= 24'b000001000000001000100110;
#10000;
	data_in <= 24'b000001100000001100101010;
#10000;
	data_in <= 24'b000001110000010100101111;
#10000;
	data_in <= 24'b000010000000011100110011;
#10000;
	data_in <= 24'b000000110000001000011100;
#10000;
	data_in <= 24'b000001000000001000011111;
#10000;
	data_in <= 24'b000001100000010000100010;
#10000;
	data_in <= 24'b000001110000001100100110;
#10000;
	data_in <= 24'b000001100000010000101000;
#10000;
	data_in <= 24'b000001110000001100101100;
#10000;
	data_in <= 24'b000010000000010100110010;
#10000;
	data_in <= 24'b000010010000011100110101;
#10000;
	data_in <= 24'b000000110000001000011100;
#10000;
	data_in <= 24'b000001010000001100100000;
#10000;
	data_in <= 24'b000001100000010000100010;
#10000;
	data_in <= 24'b000001110000001100100110;
#10000;
	data_in <= 24'b000001100000001100101010;
#10000;
	data_in <= 24'b000001110000001100101100;
#10000;
	data_in <= 24'b000001110000010000110001;
#10000;
	data_in <= 24'b000001110000010100110011;
#10000;
	data_in <= 24'b000000100000000100011011;
#10000;
	data_in <= 24'b000001000000001000011111;
#10000;
	data_in <= 24'b000001100000010000100010;
#10000;
	data_in <= 24'b000001110000001100100110;
#10000;
	data_in <= 24'b000001010000001000101001;
#10000;
	data_in <= 24'b000001010000000100101011;
#10000;
	data_in <= 24'b000001000000000100101110;
#10000;
	data_in <= 24'b000001010000001100110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001000000010100101011;
#10000;
	data_in <= 24'b000001110000011100101111;
#10000;
	data_in <= 24'b000001100000100000110001;
#10000;
	data_in <= 24'b000001000000011100110011;
#10000;
	data_in <= 24'b000001100000100100110110;
#10000;
	data_in <= 24'b000001010000100100111010;
#10000;
	data_in <= 24'b000001100000100100111100;
#10000;
	data_in <= 24'b000010100000110001000010;
#10000;
	data_in <= 24'b000001010000010100101101;
#10000;
	data_in <= 24'b000001100000100000110001;
#10000;
	data_in <= 24'b000001010000100000110100;
#10000;
	data_in <= 24'b000001110000101000110111;
#10000;
	data_in <= 24'b000010000000110000111101;
#10000;
	data_in <= 24'b000010100000110101000000;
#10000;
	data_in <= 24'b000011010000111101000101;
#10000;
	data_in <= 24'b000100000001001101001010;
#10000;
	data_in <= 24'b000010000000011100110001;
#10000;
	data_in <= 24'b000010010000101000110110;
#10000;
	data_in <= 24'b000001110000101000110111;
#10000;
	data_in <= 24'b000001110000100100111001;
#10000;
	data_in <= 24'b000001100000100100111100;
#10000;
	data_in <= 24'b000001100000100101000000;
#10000;
	data_in <= 24'b000001110000100101000011;
#10000;
	data_in <= 24'b000010000000110001000111;
#10000;
	data_in <= 24'b000001000000001100101111;
#10000;
	data_in <= 24'b000001010000010100110011;
#10000;
	data_in <= 24'b000001000000011000110110;
#10000;
	data_in <= 24'b000000110000011100111000;
#10000;
	data_in <= 24'b000001010000100000111111;
#10000;
	data_in <= 24'b000001000000100001000010;
#10000;
	data_in <= 24'b000001100000101001000101;
#10000;
	data_in <= 24'b000010000000110101001010;
#10000;
	data_in <= 24'b000001110000010100110011;
#10000;
	data_in <= 24'b000010000000100000111000;
#10000;
	data_in <= 24'b000001110000100000111010;
#10000;
	data_in <= 24'b000001100000100100111100;
#10000;
	data_in <= 24'b000010000000101001000100;
#10000;
	data_in <= 24'b000010000000110001000111;
#10000;
	data_in <= 24'b000010100000110001001100;
#10000;
	data_in <= 24'b000011000001000001010001;
#10000;
	data_in <= 24'b000010110000100000111001;
#10000;
	data_in <= 24'b000010100000101100111101;
#10000;
	data_in <= 24'b000010100000101100111110;
#10000;
	data_in <= 24'b000001110000101101000000;
#10000;
	data_in <= 24'b000010010000101101000101;
#10000;
	data_in <= 24'b000010000000101101001000;
#10000;
	data_in <= 24'b000001110000101101001100;
#10000;
	data_in <= 24'b000010010000111101010010;
#10000;
	data_in <= 24'b000001100000001100110100;
#10000;
	data_in <= 24'b000001010000011000111000;
#10000;
	data_in <= 24'b000001110000011100111101;
#10000;
	data_in <= 24'b000001100000100101000000;
#10000;
	data_in <= 24'b000010100000101101000111;
#10000;
	data_in <= 24'b000010110000111001001011;
#10000;
	data_in <= 24'b000010110000111101010000;
#10000;
	data_in <= 24'b000011100001001101011000;
#10000;
	data_in <= 24'b000010110000100000111010;
#10000;
	data_in <= 24'b000010100000101100111110;
#10000;
	data_in <= 24'b000010110000101101000001;
#10000;
	data_in <= 24'b000010010000101101000101;
#10000;
	data_in <= 24'b000011000000110101001001;
#10000;
	data_in <= 24'b000011000000111001001110;
#10000;
	data_in <= 24'b000011000001000001010001;
#10000;
	data_in <= 24'b000011100001001101011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000010000000101001000000;
#10000;
	data_in <= 24'b000010000000101101000010;
#10000;
	data_in <= 24'b000010100000110101000100;
#10000;
	data_in <= 24'b000010010000110101000111;
#10000;
	data_in <= 24'b000010110000111101001010;
#10000;
	data_in <= 24'b000011010001001001001111;
#10000;
	data_in <= 24'b000011000001001101010010;
#10000;
	data_in <= 24'b000010100001001101010011;
#10000;
	data_in <= 24'b000010100000110001000110;
#10000;
	data_in <= 24'b000010100000111001001000;
#10000;
	data_in <= 24'b000011000001000001001011;
#10000;
	data_in <= 24'b000011000001000101001110;
#10000;
	data_in <= 24'b000011100001001101010010;
#10000;
	data_in <= 24'b000011110001010101010110;
#10000;
	data_in <= 24'b000011010001010001011001;
#10000;
	data_in <= 24'b000010110001001101011001;
#10000;
	data_in <= 24'b000010100000110101001010;
#10000;
	data_in <= 24'b000010110001000001001101;
#10000;
	data_in <= 24'b000011100001001101010010;
#10000;
	data_in <= 24'b000011100001010001010101;
#10000;
	data_in <= 24'b000011110001010101011000;
#10000;
	data_in <= 24'b000011110001011001011011;
#10000;
	data_in <= 24'b000011110001011001011111;
#10000;
	data_in <= 24'b000011000001010101011111;
#10000;
	data_in <= 24'b000010010000110101001110;
#10000;
	data_in <= 24'b000010100001000001010001;
#10000;
	data_in <= 24'b000011000001001001010101;
#10000;
	data_in <= 24'b000010110001001001010111;
#10000;
	data_in <= 24'b000011010001001101011100;
#10000;
	data_in <= 24'b000011100001010001011111;
#10000;
	data_in <= 24'b000011010001010001100011;
#10000;
	data_in <= 24'b000010100001001101100011;
#10000;
	data_in <= 24'b000010010000111001010011;
#10000;
	data_in <= 24'b000010010000111101010110;
#10000;
	data_in <= 24'b000010110001000101011010;
#10000;
	data_in <= 24'b000010100001000101011010;
#10000;
	data_in <= 24'b000010110001000101011110;
#10000;
	data_in <= 24'b000011000001001101100010;
#10000;
	data_in <= 24'b000011100001010001100111;
#10000;
	data_in <= 24'b000011010001010001101001;
#10000;
	data_in <= 24'b000010100001000001011001;
#10000;
	data_in <= 24'b000011000001001001011101;
#10000;
	data_in <= 24'b000011010001001101100000;
#10000;
	data_in <= 24'b000010110001001001100001;
#10000;
	data_in <= 24'b000011000001001101100011;
#10000;
	data_in <= 24'b000011010001010001101001;
#10000;
	data_in <= 24'b000100000001011101101110;
#10000;
	data_in <= 24'b000011110001011101110001;
#10000;
	data_in <= 24'b000011000001000101011100;
#10000;
	data_in <= 24'b000011100001001101100010;
#10000;
	data_in <= 24'b000100000001010001100101;
#10000;
	data_in <= 24'b000011100001010001100111;
#10000;
	data_in <= 24'b000011110001010001101001;
#10000;
	data_in <= 24'b000100000001011001101111;
#10000;
	data_in <= 24'b000100110001100001110011;
#10000;
	data_in <= 24'b000100100001100001110111;
#10000;
	data_in <= 24'b000011000001000001011110;
#10000;
	data_in <= 24'b000011100001001101100010;
#10000;
	data_in <= 24'b000011110001010101101000;
#10000;
	data_in <= 24'b000100000001010101101010;
#10000;
	data_in <= 24'b000011110001011001101101;
#10000;
	data_in <= 24'b000100010001011001110001;
#10000;
	data_in <= 24'b000100010001100001110101;
#10000;
	data_in <= 24'b000100100001100001111001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000010010001001001010110;
#10000;
	data_in <= 24'b000010010001010001011000;
#10000;
	data_in <= 24'b000010100001011001011110;
#10000;
	data_in <= 24'b000010110001100101100001;
#10000;
	data_in <= 24'b000010110001100001100010;
#10000;
	data_in <= 24'b000010110001100101100101;
#10000;
	data_in <= 24'b000011110001110001101010;
#10000;
	data_in <= 24'b000100010010000001101111;
#10000;
	data_in <= 24'b000011110001100001100001;
#10000;
	data_in <= 24'b000011100001100101100011;
#10000;
	data_in <= 24'b000011010001101001100110;
#10000;
	data_in <= 24'b000011110001110001101010;
#10000;
	data_in <= 24'b000100000001110101101100;
#10000;
	data_in <= 24'b000011110001111001101101;
#10000;
	data_in <= 24'b000100010001111101110001;
#10000;
	data_in <= 24'b000100100010001001110101;
#10000;
	data_in <= 24'b000011100001100001100101;
#10000;
	data_in <= 24'b000010110001011101100101;
#10000;
	data_in <= 24'b000011000001011101101001;
#10000;
	data_in <= 24'b000011100001100101101101;
#10000;
	data_in <= 24'b000100000001101101101111;
#10000;
	data_in <= 24'b000011110001110001110010;
#10000;
	data_in <= 24'b000100010001110101110101;
#10000;
	data_in <= 24'b000100010001111101111000;
#10000;
	data_in <= 24'b000010010001010001100110;
#10000;
	data_in <= 24'b000010010001010001101000;
#10000;
	data_in <= 24'b000010110001010101101101;
#10000;
	data_in <= 24'b000010110001011001110000;
#10000;
	data_in <= 24'b000011010001100001110010;
#10000;
	data_in <= 24'b000011010001101001110110;
#10000;
	data_in <= 24'b000100000001110101111001;
#10000;
	data_in <= 24'b000011110001110101111101;
#10000;
	data_in <= 24'b000011010001010101101110;
#10000;
	data_in <= 24'b000011110001100001110010;
#10000;
	data_in <= 24'b000100100001101001110111;
#10000;
	data_in <= 24'b000100010001101101111001;
#10000;
	data_in <= 24'b000100010001101001111011;
#10000;
	data_in <= 24'b000100010001110001111110;
#10000;
	data_in <= 24'b000101010010000010000010;
#10000;
	data_in <= 24'b000100110010000110000111;
#10000;
	data_in <= 24'b000011100001011001110011;
#10000;
	data_in <= 24'b000100100001100101111010;
#10000;
	data_in <= 24'b000100110001110001111110;
#10000;
	data_in <= 24'b000100010001101110000000;
#10000;
	data_in <= 24'b000100000001100110000000;
#10000;
	data_in <= 24'b000100100001101110000010;
#10000;
	data_in <= 24'b000100110001111010000110;
#10000;
	data_in <= 24'b000100110010000010001010;
#10000;
	data_in <= 24'b000011110001011001110111;
#10000;
	data_in <= 24'b000100100001011101111101;
#10000;
	data_in <= 24'b000100100001100110000000;
#10000;
	data_in <= 24'b000100000001100110000001;
#10000;
	data_in <= 24'b000100000001100010000011;
#10000;
	data_in <= 24'b000100010001101110000110;
#10000;
	data_in <= 24'b000100110001110110001001;
#10000;
	data_in <= 24'b000100100001110110001100;
#10000;
	data_in <= 24'b000100110001100101111100;
#10000;
	data_in <= 24'b000100110001101010000001;
#10000;
	data_in <= 24'b000101010001101110000100;
#10000;
	data_in <= 24'b000100110001101110000110;
#10000;
	data_in <= 24'b000100110001110110001001;
#10000;
	data_in <= 24'b000101110010000110001101;
#10000;
	data_in <= 24'b000110010010001010010001;
#10000;
	data_in <= 24'b000101110010001010010001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000100010010000101110100;
#10000;
	data_in <= 24'b000100010010001001111000;
#10000;
	data_in <= 24'b000100100010000101110111;
#10000;
	data_in <= 24'b000101100010011101111110;
#10000;
	data_in <= 24'b000011100001111101110110;
#10000;
	data_in <= 24'b000010100001110101110100;
#10000;
	data_in <= 24'b000001100001100101110000;
#10000;
	data_in <= 24'b000011010001111101111000;
#10000;
	data_in <= 24'b000100100010001001111011;
#10000;
	data_in <= 24'b000010110001110101111000;
#10000;
	data_in <= 24'b000111100010110110001001;
#10000;
	data_in <= 24'b001011100100000010011011;
#10000;
	data_in <= 24'b000010010001101001110111;
#10000;
	data_in <= 24'b000011100001111101111100;
#10000;
	data_in <= 24'b000101010010011010000011;
#10000;
	data_in <= 24'b000011110010000001111101;
#10000;
	data_in <= 24'b000010100001101001111010;
#10000;
	data_in <= 24'b000100100010001110000100;
#10000;
	data_in <= 24'b001000100011001010010011;
#10000;
	data_in <= 24'b001011000011110110011110;
#10000;
	data_in <= 24'b000101110010011110001011;
#10000;
	data_in <= 24'b000100000010000010000100;
#10000;
	data_in <= 24'b000011110001111110000011;
#10000;
	data_in <= 24'b000100010010000110000101;
#10000;
	data_in <= 24'b000010100001100101111101;
#10000;
	data_in <= 24'b000101110010011010001100;
#10000;
	data_in <= 24'b000111010010110010010011;
#10000;
	data_in <= 24'b000101110010011010001101;
#10000;
	data_in <= 24'b001001010011010010011011;
#10000;
	data_in <= 24'b000100000001111110000110;
#10000;
	data_in <= 24'b000001110001011001111101;
#10000;
	data_in <= 24'b000011110001111010000101;
#10000;
	data_in <= 24'b000101000010001010001100;
#10000;
	data_in <= 24'b000011110001111110001010;
#10000;
	data_in <= 24'b000101100010011010010001;
#10000;
	data_in <= 24'b000100010010000110001100;
#10000;
	data_in <= 24'b000111000010110010010111;
#10000;
	data_in <= 24'b000011110001111110001010;
#10000;
	data_in <= 24'b000100010010000110001100;
#10000;
	data_in <= 24'b000011010001110110001000;
#10000;
	data_in <= 24'b000101110010010010010010;
#10000;
	data_in <= 24'b000011110001111010001100;
#10000;
	data_in <= 24'b000100100010000010010000;
#10000;
	data_in <= 24'b000101010010010010010010;
#10000;
	data_in <= 24'b000100010001111110001111;
#10000;
	data_in <= 24'b000100110010001010010000;
#10000;
	data_in <= 24'b000110000010011010010110;
#10000;
	data_in <= 24'b000101010010001110010011;
#10000;
	data_in <= 24'b000101010010000110010001;
#10000;
	data_in <= 24'b000101010010001110010011;
#10000;
	data_in <= 24'b000100100010000010010001;
#10000;
	data_in <= 24'b000101000010001010010010;
#10000;
	data_in <= 24'b000101000010001010010011;
#10000;
	data_in <= 24'b000101100010010010010100;
#10000;
	data_in <= 24'b000101010010001110010100;
#10000;
	data_in <= 24'b000110100010100010011001;
#10000;
	data_in <= 24'b000110000010001110010101;
#10000;
	data_in <= 24'b000100110010000110010010;
#10000;
	data_in <= 24'b000101110010010110010110;
#10000;
	data_in <= 24'b000101010010001110010100;
#10000;
	data_in <= 24'b000110100010100010011001;
#10000;
	data_in <= 24'b000101010010001110010100;
#10000;
	data_in <= 24'b000110000010011010010111;
#10000;
	data_in <= 24'b000101100010010010010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000010110001110101110110;
#10000;
	data_in <= 24'b000100000010001001111011;
#10000;
	data_in <= 24'b000101000010011001111111;
#10000;
	data_in <= 24'b000100100010010101111100;
#10000;
	data_in <= 24'b000100010010010001111011;
#10000;
	data_in <= 24'b000100010010010001111011;
#10000;
	data_in <= 24'b000100000010001101111010;
#10000;
	data_in <= 24'b000011100010000101111000;
#10000;
	data_in <= 24'b000011110010000001111101;
#10000;
	data_in <= 24'b000101000010010110000010;
#10000;
	data_in <= 24'b000101100010011110000100;
#10000;
	data_in <= 24'b000101000010010110000010;
#10000;
	data_in <= 24'b000100100010001110000000;
#10000;
	data_in <= 24'b000100110010010110000000;
#10000;
	data_in <= 24'b000100100010001110000000;
#10000;
	data_in <= 24'b000100000010001001111101;
#10000;
	data_in <= 24'b000011110001111110000011;
#10000;
	data_in <= 24'b000100100010001010000110;
#10000;
	data_in <= 24'b000100110010001110000111;
#10000;
	data_in <= 24'b000100010010000110000101;
#10000;
	data_in <= 24'b000100000010000010000100;
#10000;
	data_in <= 24'b000100010010001010000011;
#10000;
	data_in <= 24'b000100100010001010000110;
#10000;
	data_in <= 24'b000100010010001010000011;
#10000;
	data_in <= 24'b000100000001111110000110;
#10000;
	data_in <= 24'b000100010010000010000111;
#10000;
	data_in <= 24'b000100100010000110001000;
#10000;
	data_in <= 24'b000100000001111110000110;
#10000;
	data_in <= 24'b000100010010000010000111;
#10000;
	data_in <= 24'b000100110010001010001001;
#10000;
	data_in <= 24'b000101000010001110001010;
#10000;
	data_in <= 24'b000101000010001110001010;
#10000;
	data_in <= 24'b000100110010001110001110;
#10000;
	data_in <= 24'b000100110010001110001110;
#10000;
	data_in <= 24'b000100100010000110001111;
#10000;
	data_in <= 24'b000100010010000010001110;
#10000;
	data_in <= 24'b000100100010000110001111;
#10000;
	data_in <= 24'b000101000010001110010001;
#10000;
	data_in <= 24'b000101010010010010010010;
#10000;
	data_in <= 24'b000101010010010010010010;
#10000;
	data_in <= 24'b000101010010001110010011;
#10000;
	data_in <= 24'b000101000010001010010010;
#10000;
	data_in <= 24'b000100110010000110010001;
#10000;
	data_in <= 24'b000100100010000010010001;
#10000;
	data_in <= 24'b000100110010000110010010;
#10000;
	data_in <= 24'b000101000010001010010011;
#10000;
	data_in <= 24'b000100110010000110010010;
#10000;
	data_in <= 24'b000100110010000110010010;
#10000;
	data_in <= 24'b000101110010010110010110;
#10000;
	data_in <= 24'b000101010010001110010100;
#10000;
	data_in <= 24'b000101000010001010010011;
#10000;
	data_in <= 24'b000101000010000110010101;
#10000;
	data_in <= 24'b000100110010001010010110;
#10000;
	data_in <= 24'b000100100010000110010101;
#10000;
	data_in <= 24'b000100010010000010010100;
#10000;
	data_in <= 24'b000100100001111010010100;
#10000;
	data_in <= 24'b000110100010011110011011;
#10000;
	data_in <= 24'b000110010010011010011010;
#10000;
	data_in <= 24'b000110000010010110011001;
#10000;
	data_in <= 24'b000110010010011010011010;
#10000;
	data_in <= 24'b000110000010011010011100;
#10000;
	data_in <= 24'b000110000010011010011100;
#10000;
	data_in <= 24'b000101100010010010011010;
#10000;
	data_in <= 24'b000101000010001010011000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000011110010000001110111;
#10000;
	data_in <= 24'b000101000010010101111011;
#10000;
	data_in <= 24'b000101010010011001111100;
#10000;
	data_in <= 24'b000100010010000101110100;
#10000;
	data_in <= 24'b000011110001110101101111;
#10000;
	data_in <= 24'b000100000001110101101100;
#10000;
	data_in <= 24'b000011010001101001101001;
#10000;
	data_in <= 24'b000010100001011101100011;
#10000;
	data_in <= 24'b000101000010001101111111;
#10000;
	data_in <= 24'b000100110010001001111110;
#10000;
	data_in <= 24'b000100000001111101111011;
#10000;
	data_in <= 24'b000011100001111001110111;
#10000;
	data_in <= 24'b000011110001110101110101;
#10000;
	data_in <= 24'b000100010001111001110100;
#10000;
	data_in <= 24'b000100000001111001110001;
#10000;
	data_in <= 24'b000100100001111001110000;
#10000;
	data_in <= 24'b000100100010001010000011;
#10000;
	data_in <= 24'b000011100001111001111110;
#10000;
	data_in <= 24'b000011000001110001111100;
#10000;
	data_in <= 24'b000100010010000001111101;
#10000;
	data_in <= 24'b000100110010001001111111;
#10000;
	data_in <= 24'b000100100001111101111011;
#10000;
	data_in <= 24'b000011110001110101110110;
#10000;
	data_in <= 24'b000100000001110001110100;
#10000;
	data_in <= 24'b000101000010000110001001;
#10000;
	data_in <= 24'b000100100010000010000110;
#10000;
	data_in <= 24'b000100010001111110000101;
#10000;
	data_in <= 24'b000100100010000110000101;
#10000;
	data_in <= 24'b000101010010000110000110;
#10000;
	data_in <= 24'b000100110010000010000010;
#10000;
	data_in <= 24'b000100000001110001111100;
#10000;
	data_in <= 24'b000011010001100101110111;
#10000;
	data_in <= 24'b000110010010011010010100;
#10000;
	data_in <= 24'b000110010010011010010100;
#10000;
	data_in <= 24'b000101010010001010010000;
#10000;
	data_in <= 24'b000100000001110110001001;
#10000;
	data_in <= 24'b000100000001110110000111;
#10000;
	data_in <= 24'b000100100001111110000111;
#10000;
	data_in <= 24'b000100110001111110000101;
#10000;
	data_in <= 24'b000100000001110010000001;
#10000;
	data_in <= 24'b000101010001111110010100;
#10000;
	data_in <= 24'b000110010010001110011000;
#10000;
	data_in <= 24'b000110000010001110010101;
#10000;
	data_in <= 24'b000100110001111010010000;
#10000;
	data_in <= 24'b000100100001110110001101;
#10000;
	data_in <= 24'b000101010010000010001111;
#10000;
	data_in <= 24'b000101110010000110001101;
#10000;
	data_in <= 24'b000100110001111010000110;
#10000;
	data_in <= 24'b000100100001101110010100;
#10000;
	data_in <= 24'b000101010001111010010111;
#10000;
	data_in <= 24'b000101100001111110011000;
#10000;
	data_in <= 24'b000101100010000010010110;
#10000;
	data_in <= 24'b000101100010000010010101;
#10000;
	data_in <= 24'b000101110010001010010100;
#10000;
	data_in <= 24'b000101100010000110010001;
#10000;
	data_in <= 24'b000101000010000010001100;
#10000;
	data_in <= 24'b000101110001111110011010;
#10000;
	data_in <= 24'b000101010001110110011000;
#10000;
	data_in <= 24'b000101000001110010010111;
#10000;
	data_in <= 24'b000101010001111010010111;
#10000;
	data_in <= 24'b000101110010000010011001;
#10000;
	data_in <= 24'b000101110010000110010110;
#10000;
	data_in <= 24'b000110100010010010010110;
#10000;
	data_in <= 24'b000110110010011010010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000011100001100101100011;
#10000;
	data_in <= 24'b000011110001100001100001;
#10000;
	data_in <= 24'b000011000001011001011100;
#10000;
	data_in <= 24'b000011000001010101011001;
#10000;
	data_in <= 24'b000011010001010101011000;
#10000;
	data_in <= 24'b000100000001011001011001;
#10000;
	data_in <= 24'b000011110001010101010110;
#10000;
	data_in <= 24'b000011100001010101010100;
#10000;
	data_in <= 24'b000100110001111001101110;
#10000;
	data_in <= 24'b000101000001111001101100;
#10000;
	data_in <= 24'b000100100001110101100111;
#10000;
	data_in <= 24'b000100100001101101100100;
#10000;
	data_in <= 24'b000100110001101001100011;
#10000;
	data_in <= 24'b000100100001101001100000;
#10000;
	data_in <= 24'b000100000001100001011110;
#10000;
	data_in <= 24'b000011010001011001011001;
#10000;
	data_in <= 24'b000011010001100001101100;
#10000;
	data_in <= 24'b000011100001100101101011;
#10000;
	data_in <= 24'b000011010001100001101000;
#10000;
	data_in <= 24'b000011100001100001100110;
#10000;
	data_in <= 24'b000011110001100101100110;
#10000;
	data_in <= 24'b000100110001110001100110;
#10000;
	data_in <= 24'b000100110001110001100110;
#10000;
	data_in <= 24'b000100010001101001100011;
#10000;
	data_in <= 24'b000011110001101001110100;
#10000;
	data_in <= 24'b000011010001100101110001;
#10000;
	data_in <= 24'b000010110001010101101100;
#10000;
	data_in <= 24'b000010000001001101100111;
#10000;
	data_in <= 24'b000010100001010101100111;
#10000;
	data_in <= 24'b000011000001011101100111;
#10000;
	data_in <= 24'b000010110001011001100110;
#10000;
	data_in <= 24'b000010100001011001100100;
#10000;
	data_in <= 24'b000100000001110001111100;
#10000;
	data_in <= 24'b000011110001101101111001;
#10000;
	data_in <= 24'b000011100001100101110101;
#10000;
	data_in <= 24'b000011000001011101110001;
#10000;
	data_in <= 24'b000011110001100101110001;
#10000;
	data_in <= 24'b000100000001101001110001;
#10000;
	data_in <= 24'b000011100001100001101111;
#10000;
	data_in <= 24'b000010110001011001101010;
#10000;
	data_in <= 24'b000011100001101010000000;
#10000;
	data_in <= 24'b000011100001101001111111;
#10000;
	data_in <= 24'b000100000001101101111101;
#10000;
	data_in <= 24'b000100010001110101111101;
#10000;
	data_in <= 24'b000100110001111101111101;
#10000;
	data_in <= 24'b000101000010000101111101;
#10000;
	data_in <= 24'b000100110001111001111010;
#10000;
	data_in <= 24'b000011110001101101110011;
#10000;
	data_in <= 24'b000100110010000010001010;
#10000;
	data_in <= 24'b000100100001111110000111;
#10000;
	data_in <= 24'b000100100001111010000100;
#10000;
	data_in <= 24'b000100100001111010000011;
#10000;
	data_in <= 24'b000100110010000010000010;
#10000;
	data_in <= 24'b000100100010000010000000;
#10000;
	data_in <= 24'b000100010001110101111101;
#10000;
	data_in <= 24'b000011000001100001110110;
#10000;
	data_in <= 24'b000101010010000010001111;
#10000;
	data_in <= 24'b000100110010000010001010;
#10000;
	data_in <= 24'b000100100001110110000101;
#10000;
	data_in <= 24'b000100010001110110000011;
#10000;
	data_in <= 24'b000101000010000010000101;
#10000;
	data_in <= 24'b000101110010001110001000;
#10000;
	data_in <= 24'b000101110010010010000110;
#10000;
	data_in <= 24'b000101000010001010000010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000011110001011101010011;
#10000;
	data_in <= 24'b000011010001010101010000;
#10000;
	data_in <= 24'b000010110001001101001110;
#10000;
	data_in <= 24'b000011000001001101001100;
#10000;
	data_in <= 24'b000011010001001001001001;
#10000;
	data_in <= 24'b000010100001000101000011;
#10000;
	data_in <= 24'b000010010000111000111111;
#10000;
	data_in <= 24'b000001110000101100111011;
#10000;
	data_in <= 24'b000010010001001101010011;
#10000;
	data_in <= 24'b000010110001010001010011;
#10000;
	data_in <= 24'b000011000001010101010100;
#10000;
	data_in <= 24'b000011000001010001010000;
#10000;
	data_in <= 24'b000010110001000101001100;
#10000;
	data_in <= 24'b000010110001000001000111;
#10000;
	data_in <= 24'b000010110001000101000110;
#10000;
	data_in <= 24'b000011010001001001000011;
#10000;
	data_in <= 24'b000011010001011101011101;
#10000;
	data_in <= 24'b000011010001100101011011;
#10000;
	data_in <= 24'b000011100001011101011010;
#10000;
	data_in <= 24'b000011000001010101010101;
#10000;
	data_in <= 24'b000010100001000101010000;
#10000;
	data_in <= 24'b000010010000111101001010;
#10000;
	data_in <= 24'b000010010000110101000111;
#10000;
	data_in <= 24'b000010100000111001000011;
#10000;
	data_in <= 24'b000010100001011101100001;
#10000;
	data_in <= 24'b000010010001010101011101;
#10000;
	data_in <= 24'b000010010001001001011011;
#10000;
	data_in <= 24'b000010110001010001011000;
#10000;
	data_in <= 24'b000011100001011001011001;
#10000;
	data_in <= 24'b000100010001100001010111;
#10000;
	data_in <= 24'b000011110001010001010001;
#10000;
	data_in <= 24'b000011000001000001001010;
#10000;
	data_in <= 24'b000011010001101001101001;
#10000;
	data_in <= 24'b000011000001100001100110;
#10000;
	data_in <= 24'b000011000001011001100011;
#10000;
	data_in <= 24'b000011010001011001100000;
#10000;
	data_in <= 24'b000100010001100001100001;
#10000;
	data_in <= 24'b000100100001100101011110;
#10000;
	data_in <= 24'b000100010001010001011000;
#10000;
	data_in <= 24'b000011010000111101001111;
#10000;
	data_in <= 24'b000100000001110101110011;
#10000;
	data_in <= 24'b000100110001111101110001;
#10000;
	data_in <= 24'b000100100001110101101111;
#10000;
	data_in <= 24'b000011110001100101100111;
#10000;
	data_in <= 24'b000011000001010001100001;
#10000;
	data_in <= 24'b000010110001001001011011;
#10000;
	data_in <= 24'b000010110000111101010110;
#10000;
	data_in <= 24'b000010100000110101010001;
#10000;
	data_in <= 24'b000011110001101001110100;
#10000;
	data_in <= 24'b000100100001110001110011;
#10000;
	data_in <= 24'b000100100001101101110010;
#10000;
	data_in <= 24'b000011100001011001101001;
#10000;
	data_in <= 24'b000010110001001001100010;
#10000;
	data_in <= 24'b000011010001001101100000;
#10000;
	data_in <= 24'b000100010001010001011111;
#10000;
	data_in <= 24'b000100100001010001011011;
#10000;
	data_in <= 24'b000110000010001101111111;
#10000;
	data_in <= 24'b000101100010001001111010;
#10000;
	data_in <= 24'b000100110001101101110100;
#10000;
	data_in <= 24'b000011000001011001101010;
#10000;
	data_in <= 24'b000011100001010001100111;
#10000;
	data_in <= 24'b000100100001011101100110;
#10000;
	data_in <= 24'b000100100001011001100100;
#10000;
	data_in <= 24'b000100010001010001011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001110000101000110110;
#10000;
	data_in <= 24'b000010110000111100111000;
#10000;
	data_in <= 24'b000010110001000000110111;
#10000;
	data_in <= 24'b000010100001000000110101;
#10000;
	data_in <= 24'b000010110000111000110100;
#10000;
	data_in <= 24'b000010000000101100110001;
#10000;
	data_in <= 24'b000001100000100100101111;
#10000;
	data_in <= 24'b000001100000101000101101;
#10000;
	data_in <= 24'b000001110000101100111011;
#10000;
	data_in <= 24'b000010100000110100111001;
#10000;
	data_in <= 24'b000010010000110000111000;
#10000;
	data_in <= 24'b000010010000110100110110;
#10000;
	data_in <= 24'b000011000001000100111000;
#10000;
	data_in <= 24'b000010100000111100110110;
#10000;
	data_in <= 24'b000001110000100100110001;
#10000;
	data_in <= 24'b000001100000100000110000;
#10000;
	data_in <= 24'b000100000001001101000110;
#10000;
	data_in <= 24'b000011010001000101000001;
#10000;
	data_in <= 24'b000010010000110100111101;
#10000;
	data_in <= 24'b000010010000111000111011;
#10000;
	data_in <= 24'b000011010001001100111110;
#10000;
	data_in <= 24'b000011000001001000111011;
#10000;
	data_in <= 24'b000010000000110000110101;
#10000;
	data_in <= 24'b000001100000101000110011;
#10000;
	data_in <= 24'b000101110001101001010001;
#10000;
	data_in <= 24'b000100110001010101001011;
#10000;
	data_in <= 24'b000011000000111101000010;
#10000;
	data_in <= 24'b000010100000111000111110;
#10000;
	data_in <= 24'b000011010001000101000001;
#10000;
	data_in <= 24'b000011000001000100111110;
#10000;
	data_in <= 24'b000010000000111000111001;
#10000;
	data_in <= 24'b000001110000110100111000;
#10000;
	data_in <= 24'b000100110001010001010001;
#10000;
	data_in <= 24'b000100000001001001001100;
#10000;
	data_in <= 24'b000010110000111001000101;
#10000;
	data_in <= 24'b000010100000111001000001;
#10000;
	data_in <= 24'b000011000001000001000011;
#10000;
	data_in <= 24'b000010100000111101000000;
#10000;
	data_in <= 24'b000010000000110100111110;
#10000;
	data_in <= 24'b000010100000111000111111;
#10000;
	data_in <= 24'b000010010000101101001100;
#10000;
	data_in <= 24'b000011000000110101001010;
#10000;
	data_in <= 24'b000011000000110101001001;
#10000;
	data_in <= 24'b000011100001000101001000;
#10000;
	data_in <= 24'b000011110001001001001001;
#10000;
	data_in <= 24'b000010110000111101000100;
#10000;
	data_in <= 24'b000010100000111001000011;
#10000;
	data_in <= 24'b000011100001001001000111;
#10000;
	data_in <= 24'b000010110000110001010000;
#10000;
	data_in <= 24'b000011010000111101010000;
#10000;
	data_in <= 24'b000011110000111101001111;
#10000;
	data_in <= 24'b000100000001000101001101;
#10000;
	data_in <= 24'b000100000001000101001101;
#10000;
	data_in <= 24'b000011000000111001001000;
#10000;
	data_in <= 24'b000010100000111101000110;
#10000;
	data_in <= 24'b000100010001010001001011;
#10000;
	data_in <= 24'b000100110001001101011001;
#10000;
	data_in <= 24'b000100100001010001010101;
#10000;
	data_in <= 24'b000100010001000001010010;
#10000;
	data_in <= 24'b000011110001000001001101;
#10000;
	data_in <= 24'b000011010000111001001011;
#10000;
	data_in <= 24'b000010100000101101000111;
#10000;
	data_in <= 24'b000010010000110101000111;
#10000;
	data_in <= 24'b000100000001010001001110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
	data_in <= 24'b000001010000100100101100;
#10000;
	data_in <= 24'b000001000000100000101011;
#10000;
	data_in <= 24'b000010010000111000101111;
#10000;
	data_in <= 24'b000011000001000100110010;
#10000;
	data_in <= 24'b000011110001000100110011;
#10000;
	data_in <= 24'b000010110000111000101101;
#10000;
	data_in <= 24'b000001000000011100100110;
#10000;
	data_in <= 24'b000010010000110000101011;
#10000;
	data_in <= 24'b000011000000111000110110;
#10000;
	data_in <= 24'b000010010000101100110011;
#10000;
	data_in <= 24'b000010010000110000110010;
#10000;
	data_in <= 24'b000001100000100100101111;
#10000;
	data_in <= 24'b000010000000101000101101;
#10000;
	data_in <= 24'b000001110000100100101100;
#10000;
	data_in <= 24'b000001010000011100101010;
#10000;
	data_in <= 24'b000011010000111100110001;
#10000;
	data_in <= 24'b000001110000101100110100;
#10000;
	data_in <= 24'b000010000000110000110101;
#10000;
	data_in <= 24'b000010110000110100110110;
#10000;
	data_in <= 24'b000001110000100100110010;
#10000;
	data_in <= 24'b000001110000100100110001;
#10000;
	data_in <= 24'b000010000000101000110010;
#10000;
	data_in <= 24'b000001010000100000101110;
#10000;
	data_in <= 24'b000010100000110100110011;
#10000;
	data_in <= 24'b000001010000100000110101;
#10000;
	data_in <= 24'b000010010000110000111001;
#10000;
	data_in <= 24'b000011100000111000111100;
#10000;
	data_in <= 24'b000010100000101100110111;
#10000;
	data_in <= 24'b000010100000101100110111;
#10000;
	data_in <= 24'b000010100000110000110101;
#10000;
	data_in <= 24'b000001100000100000110001;
#10000;
	data_in <= 24'b000010000000101000110010;
#10000;
	data_in <= 24'b000011110001000001000010;
#10000;
	data_in <= 24'b000011110001000001000010;
#10000;
	data_in <= 24'b000011100001000001000000;
#10000;
	data_in <= 24'b000001100000100000111000;
#10000;
	data_in <= 24'b000001010000011100110111;
#10000;
	data_in <= 24'b000001110000101000110111;
#10000;
	data_in <= 24'b000001100000011000110100;
#10000;
	data_in <= 24'b000010000000100100110101;
#10000;
	data_in <= 24'b000011110001000101000111;
#10000;
	data_in <= 24'b000100000001000101000100;
#10000;
	data_in <= 24'b000011100000111101000010;
#10000;
	data_in <= 24'b000001110000100000111010;
#10000;
	data_in <= 24'b000001110000100000111010;
#10000;
	data_in <= 24'b000010100000110000111100;
#10000;
	data_in <= 24'b000010000000100000111000;
#10000;
	data_in <= 24'b000010100000101000111000;
#10000;
	data_in <= 24'b000011000000110101000101;
#10000;
	data_in <= 24'b000010110000110101000011;
#10000;
	data_in <= 24'b000011100000111001000100;
#10000;
	data_in <= 24'b000010110000110000111111;
#10000;
	data_in <= 24'b000011100000111101000010;
#10000;
	data_in <= 24'b000011110001000001000010;
#10000;
	data_in <= 24'b000010100000100100111011;
#10000;
	data_in <= 24'b000010110000101100111011;
#10000;
	data_in <= 24'b000100000001000101001001;
#10000;
	data_in <= 24'b000011010000111001000110;
#10000;
	data_in <= 24'b000011100000111001000100;
#10000;
	data_in <= 24'b000011000000110001000010;
#10000;
	data_in <= 24'b000011110001000001000011;
#10000;
	data_in <= 24'b000011110001000001000011;
#10000;
	data_in <= 24'b000010100000100100111011;
#10000;
	data_in <= 24'b000010110000101100111011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
end_of_file_signal  <= 1'b1;
	data_in <= 24'b000010110000110100101100;
#10000;
	data_in <= 24'b000001100000100000100110;
#10000;
	data_in <= 24'b000001110000100100100111;
#10000;
	data_in <= 24'b000001110000101000100110;
#10000;
	data_in <= 24'b000001100000100100100101;
#10000;
	data_in <= 24'b000001000000100000100001;
#10000;
	data_in <= 24'b000000000000001100011111;
#10000;
	data_in <= 24'b000000100000011000011111;
#10000;
	data_in <= 24'b000010100000101100101101;
#10000;
	data_in <= 24'b000001010000011100100110;
#10000;
	data_in <= 24'b000001010000011100100110;
#10000;
	data_in <= 24'b000001010000011100100101;
#10000;
	data_in <= 24'b000001010000011100100101;
#10000;
	data_in <= 24'b000001100000100100100101;
#10000;
	data_in <= 24'b000001000000011000100100;
#10000;
	data_in <= 24'b000010000000101100100111;
#10000;
	data_in <= 24'b000011000000111000110001;
#10000;
	data_in <= 24'b000001100000100000101010;
#10000;
	data_in <= 24'b000010000000100100101011;
#10000;
	data_in <= 24'b000001100000100000100111;
#10000;
	data_in <= 24'b000001010000011100100110;
#10000;
	data_in <= 24'b000001010000011100100101;
#10000;
	data_in <= 24'b000000110000010100100100;
#10000;
	data_in <= 24'b000001100000100000100110;
#10000;
	data_in <= 24'b000011000000110100110011;
#10000;
	data_in <= 24'b000010010000101100101110;
#10000;
	data_in <= 24'b000010110000101100101111;
#10000;
	data_in <= 24'b000010000000100100101011;
#10000;
	data_in <= 24'b000001100000011100101001;
#10000;
	data_in <= 24'b000001010000011000101000;
#10000;
	data_in <= 24'b000000000000000100100011;
#10000;
	data_in <= 24'b000000100000010000100011;
#10000;
	data_in <= 24'b000010010000100000110010;
#10000;
	data_in <= 24'b000001110000011100101111;
#10000;
	data_in <= 24'b000010010000100100110001;
#10000;
	data_in <= 24'b000001110000100000101110;
#10000;
	data_in <= 24'b000001110000011000101101;
#10000;
	data_in <= 24'b000001110000011100101011;
#10000;
	data_in <= 24'b000000110000001100100111;
#10000;
	data_in <= 24'b000001100000011100101001;
#10000;
	data_in <= 24'b000010100000100100110101;
#10000;
	data_in <= 24'b000010000000011100110001;
#10000;
	data_in <= 24'b000010010000100000110010;
#10000;
	data_in <= 24'b000001100000011000101110;
#10000;
	data_in <= 24'b000001100000010100101101;
#10000;
	data_in <= 24'b000010000000011100101110;
#10000;
	data_in <= 24'b000001100000010100101100;
#10000;
	data_in <= 24'b000010100000101000101110;
#10000;
	data_in <= 24'b000010100000101000111000;
#10000;
	data_in <= 24'b000010000000100100110101;
#10000;
	data_in <= 24'b000010110000101000110100;
#10000;
	data_in <= 24'b000001110000011100101111;
#10000;
	data_in <= 24'b000001100000010100101101;
#10000;
	data_in <= 24'b000010000000011100101110;
#10000;
	data_in <= 24'b000001110000011000101101;
#10000;
	data_in <= 24'b000010100000100100110000;
#10000;
	data_in <= 24'b000001110000011100110111;
#10000;
	data_in <= 24'b000001100000011100110011;
#10000;
	data_in <= 24'b000011000000101100110111;
#10000;
	data_in <= 24'b000010010000100000110010;
#10000;
	data_in <= 24'b000010010000100000110000;
#10000;
	data_in <= 24'b000010110000101000110010;
#10000;
	data_in <= 24'b000010000000011100101110;
#10000;
	data_in <= 24'b000010100000100100110000;




#10000;
#130000;
enable <= 1'b0;

#2000000; 

$finish;
end // end of stimulus process
	
always
begin : CLOCK_clk
	//this process was generated based on formula: 0 0 ns, 1 5 ns -r 10 ns
	//#<time to next event>; // <current time>
	clk = 1'b0;
	#5000; //0
	clk = 1'b1;
	#5000; //5000
end

always 	@(JPEG_bitstream or data_ready)
begin : JPEG
		if (data_ready==1'b1) 		
					$display("%h", JPEG_bitstream);						
end	


endmodule